netcdf tas_Amon_exAA02_historical_r1i1p1_195001-195012_box {
dimensions:
	lon = 20 ;
	bnds = 2 ;
	lat = 20 ;
	time = UNLIMITED ; // (4 currently)
variables:
	double lon(lon) ;
		lon:standard_name = "longitude" ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:axis = "X" ;
		lon:bounds = "lon_bnds" ;
	double lon_bnds(lon, bnds) ;
	double lat(lat) ;
		lat:standard_name = "latitude" ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:axis = "Y" ;
		lat:bounds = "lat_bnds" ;
	double lat_bnds(lat, bnds) ;
	double height ;
		height:standard_name = "height" ;
		height:long_name = "height" ;
		height:units = "m" ;
		height:positive = "up" ;
		height:axis = "Z" ;
	double time(time) ;
		time:standard_name = "time" ;
		time:long_name = "time" ;
		time:bounds = "time_bnds" ;
		time:units = "days since 1950-1-1 00:00:00" ;
		time:calendar = "standard" ;
		time:axis = "T" ;
	double time_bnds(time, bnds) ;
	float tas(time, lat, lon) ;
		tas:standard_name = "air_temperature" ;
		tas:long_name = "Near-Surface Air Temperature" ;
		tas:units = "K" ;
		tas:grid_type = "gaussian" ;
		tas:coordinates = "height" ;
		tas:_FillValue = 1.e+20f ;
		tas:missing_value = 1.e+20f ;
		tas:original_name = "T2" ;
		tas:cell_methods = "time: mean" ;
		tas:history = "2011-04-22T07:31:59Z altered by CMOR: Treated scalar dimension: \'height\'. 2011-04-22T07:31:59Z altered by CMOR: replaced missing value flag (-999) with standard missing value (1e+20). 2011-04-22T07:31:59Z altered by CMOR: Inverted axis: lat." ;
		tas:associated_files = "baseURL: http://cmip-pcmdi.llnl.gov/CMIP5/dataLocation gridspecFile: gridspec_atmos_fx_MIROC4h_historical_r0i0p0.nc areacella: areacella_fx_MIROC4h_historical_r0i0p0.nc" ;

// global attributes:
		:CDI = "Climate Data Interface version ?? (http://mpimet.mpg.de/cdi)" ;
		:Conventions = "CF-1.4" ;
		:history = "reset by cdo to create anonymous sample file" ;
		:source = "201707_compliance_checker_evaluation/work/p1.py" ;
		:institution = "CEDA" ;
		:institute_id = "CEDA" ;
		:experiment_id = "historical" ;
		:model_id = "exAA02" ;
		:forcing = "GHG, SA, Oz, LU, Sl, Vl, SS, Ds, BC, MD, OC (GHG includes CO2, N2O, methane, and fluorocarbons; Oz includes OH and H2O2)" ;
		:parent_experiment_id = "piControl" ;
		:parent_experiment_rip = "r1i1p1" ;
		:branch_time = 14600. ;
		:contact = "none" ;
		:references = "Sakamoto et al., 2011: MIROC4h -- a new high-resolution atmosphere-ocean coupled general circulation model. (in preparation); Tatebe et al., 2011: (in preparation)" ;
		:initialization_method = 1 ;
		:physics_version = 1 ;
		:tracking_id = "d7e7f8f2-f746-451c-b373-1acd1f2272b1" ;
		:product = "output" ;
		:experiment = "historical" ;
		:frequency = "mon" ;
		:creation_date = "2011-04-22T07:31:59Z" ;
		:project_id = "CMIP5" ;
		:table_id = "Table Amon (11 April 2011) 1cfdc7322cf2f4a32614826fab42c1ab" ;
		:title = "Dummy file with known metadata errors" ;
		:parent_experiment = "pre-industrial control" ;
		:modeling_realm = "atmos" ;
		:realization = 1 ;
		:cmor_version = "2.5.8" ;
		:comment = "this is a sample file with known metadata errors" ;
		:CDO = "Climate Data Operators version 1.7.0 (http://mpimet.mpg.de/cdo)" ;
data:

 lon = 0, 0.5625, 1.125, 1.6875, 2.25, 2.8125, 3.375, 3.9375, 4.5, 5.0625, 
    5.625, 6.1875, 6.75, 7.3125, 7.875, 8.4375, 9, 9.5625, 10.125, 10.6875 ;

 lon_bnds =
  -0.28125, 0.28125,
  0.28125, 0.84375,
  0.84375, 1.40625,
  1.40625, 1.96875,
  1.96875, 2.53125,
  2.53125, 3.09375,
  3.09375, 3.65625,
  3.65625, 4.21875,
  4.21875, 4.78125,
  4.78125, 5.34375,
  5.34375, 5.90625,
  5.90625, 6.46875,
  6.46875, 7.03125,
  7.03125, 7.59375,
  7.59375, 8.15625,
  8.15625, 8.71875,
  8.71875, 9.28125,
  9.28125, 9.84375,
  9.84375, 10.40625,
  10.40625, 10.96875 ;

 lat = -89.5700895506067, -89.0131761310221, -88.4529738367131, 
    -87.8920284453444, -87.3308011797376, -86.7694375145276, 
    -86.2079976214231, -85.6465108479529, -85.0849932009119, 
    -84.5234541489144, -83.9618996497181, -83.400333638737, 
    -82.8387588197095, -82.2771771114338, -81.7155899132665, 
    -81.153998269713, -80.5924029761778, -80.0308046490315, 
    -79.4692037732917, -78.907600735838 ;

 lat_bnds =
  -90, -89.3112934231673,
  -89.3112934231673, -88.7436418237873,
  -88.7436418237873, -88.1797555341309,
  -88.1797555341309, -87.6169431617971,
  -87.6169431617971, -87.054586265917,
  -87.054586265917, -86.4924650679895,
  -86.4924650679895, -85.9304816687214,
  -85.9304816687214, -85.3685858166392,
  -85.3685858166392, -84.8067490548906,
  -84.8067490548906, -84.2449540578723,
  -84.2449540578723, -83.6831896720038,
  -83.6831896720038, -83.1214483914835,
  -83.1214483914835, -82.5597249794501,
  -82.5597249794501, -81.9980156707204,
  -81.9980156707204, -81.4363176886757,
  -81.4363176886757, -80.8746289407599,
  -80.8746289407599, -80.3129478200131,
  -80.3129478200131, -79.7512730719198,
  -79.7512730719198, -79.1896037027966,
  -79.1896037027966, -78.6279389153457 ;

 height = 2 ;

 time = 15.5, 45, 74.5, 105 ;

 time_bnds =
  0, 31,
  31, 59,
  59, 90,
  90, 120 ;

 tas =
  253.4909, 253.4909, 253.4909, 253.4909, 253.4557, 253.4557, 253.4557, 
    253.4557, 253.4557, 253.4557, 253.4557, 253.4557, 253.4206, 253.4206, 
    253.4206, 253.4206, 253.4206, 253.4206, 253.4206, 253.4206,
  253.7366, 253.7366, 253.7015, 253.7015, 253.7015, 253.6664, 253.6664, 
    253.6664, 253.6313, 253.6313, 253.6313, 253.5962, 253.5962, 253.5962, 
    253.5611, 253.5611, 253.5611, 253.526, 253.526, 253.526,
  253.9473, 253.9122, 253.9122, 253.8771, 253.8419, 253.8419, 253.8068, 
    253.8068, 253.7717, 253.7366, 253.7366, 253.7015, 253.6664, 253.6313, 
    253.6313, 253.5962, 253.5611, 253.5611, 253.526, 253.4909,
  253.9473, 253.9473, 253.9122, 253.8771, 253.8419, 253.8068, 253.7717, 
    253.7717, 253.7366, 253.7015, 253.6664, 253.6313, 253.5962, 253.5611, 
    253.5611, 253.526, 253.4909, 253.4557, 253.4557, 253.4206,
  253.9824, 253.9473, 253.9122, 253.8771, 253.8771, 253.8419, 253.8068, 
    253.8068, 253.7717, 253.7366, 253.7366, 253.7015, 253.7015, 253.6664, 
    253.6664, 253.6313, 253.6313, 253.5962, 253.5962, 253.5611,
  254.0877, 254.0526, 254.0526, 254.0526, 254.0175, 254.0175, 253.9824, 
    253.9824, 253.9473, 253.9473, 253.9473, 253.9122, 253.9122, 253.8771, 
    253.8771, 253.8419, 253.8419, 253.8419, 253.8068, 253.8068,
  254.0877, 254.0877, 254.0877, 254.0526, 254.0526, 254.0526, 254.0526, 
    254.0526, 254.0175, 254.0175, 253.9824, 253.9824, 253.9473, 253.9473, 
    253.9122, 253.9122, 253.8771, 253.8771, 253.8419, 253.8068,
  253.9122, 253.9122, 253.9122, 253.9122, 253.9122, 253.9122, 253.8771, 
    253.8771, 253.8419, 253.8068, 253.8068, 253.7717, 253.7366, 253.7015, 
    253.7015, 253.6664, 253.6313, 253.5962, 253.5611, 253.526,
  253.9122, 253.9122, 253.9122, 253.9473, 253.9122, 253.9122, 253.8771, 
    253.8771, 253.8419, 253.8068, 253.8068, 253.7717, 253.7015, 253.6664, 
    253.6313, 253.5962, 253.526, 253.4909, 253.4206, 253.3504,
  254.0175, 254.0526, 254.0526, 254.0877, 254.0877, 254.0526, 254.0526, 
    254.0175, 253.9824, 253.9473, 253.9122, 253.8771, 253.8068, 253.7717, 
    253.7015, 253.6313, 253.5611, 253.4909, 253.3855, 253.3153,
  254.0877, 254.1228, 254.1228, 254.1579, 254.1579, 254.1579, 254.1228, 
    254.0877, 254.0526, 254.0175, 253.9824, 253.9122, 253.8419, 253.7717, 
    253.6664, 253.5962, 253.4909, 253.3855, 253.2802, 253.1749,
  254.1579, 254.1579, 254.1931, 254.1579, 254.1579, 254.1228, 254.0877, 
    254.0526, 253.9824, 253.9122, 253.8068, 253.7366, 253.6313, 253.526, 
    253.4206, 253.3153, 253.21, 253.0695, 252.9642, 252.8238,
  254.1931, 254.1931, 254.1931, 254.1579, 254.0877, 254.0175, 253.9473, 
    253.8771, 253.7717, 253.6664, 253.5611, 253.4206, 253.3153, 253.21, 
    253.0695, 252.9291, 252.7887, 252.6482, 252.5078, 252.4024,
  254.1579, 254.1228, 254.0877, 254.0175, 253.9473, 253.8771, 253.7717, 
    253.6664, 253.526, 253.3855, 253.2451, 253.1046, 252.9642, 252.7887, 
    252.6482, 252.5078, 252.3322, 252.1918, 252.0865, 251.9109,
  254.0175, 253.9824, 253.9122, 253.8419, 253.7717, 253.6664, 253.5611, 
    253.4206, 253.2802, 253.1046, 252.9642, 252.7887, 252.6131, 252.4375, 
    252.262, 252.0865, 251.9109, 251.7354, 251.5598, 251.4545,
  253.8771, 253.8419, 253.8068, 253.7366, 253.6313, 253.526, 253.3855, 
    253.2451, 253.0695, 252.894, 252.6833, 252.4727, 252.2971, 252.0865, 
    251.9109, 251.7354, 251.5247, 251.3842, 251.2087, 251.0683,
  253.9122, 253.8419, 253.7717, 253.7015, 253.5962, 253.4909, 253.3504, 
    253.1749, 252.9642, 252.7887, 252.578, 252.3673, 252.1216, 251.9109, 
    251.7002, 251.5247, 251.314, 251.1385, 250.9629, 250.8225,
  253.7366, 253.7015, 253.6313, 253.526, 253.4206, 253.2802, 253.1398, 
    252.9291, 252.7535, 252.5429, 252.3322, 252.0865, 251.8407, 251.63, 
    251.4194, 251.2087, 251.0332, 250.8576, 250.6821, 250.5416,
  253.4909, 253.4557, 253.3855, 253.2451, 253.1398, 252.9993, 252.8238, 
    252.6482, 252.4375, 252.1918, 251.946, 251.7002, 251.4545, 251.2087, 
    250.998, 250.8225, 250.6469, 250.5065, 250.4012, 250.2958,
  253.2451, 253.1749, 253.0344, 252.9291, 252.7887, 252.6131, 252.4024, 
    252.2269, 252.0162, 251.8056, 251.5598, 251.314, 251.0683, 250.8576, 
    250.6821, 250.5065, 250.3661, 250.2607, 250.1554, 250.0501,
  239.483, 239.483, 239.483, 239.483, 239.483, 239.444, 239.444, 239.444, 
    239.444, 239.444, 239.444, 239.444, 239.4049, 239.4049, 239.4049, 
    239.4049, 239.4049, 239.4049, 239.4049, 239.4049,
  240.1085, 240.0694, 240.0694, 240.0694, 240.0303, 240.0303, 240.0303, 
    239.9912, 239.9912, 239.9521, 239.9521, 239.9521, 239.9131, 239.9131, 
    239.9131, 239.874, 239.874, 239.874, 239.8349, 239.8349,
  240.4212, 240.3822, 240.3822, 240.3431, 240.304, 240.2649, 240.2649, 
    240.2258, 240.1867, 240.1476, 240.1476, 240.1085, 240.0694, 240.0694, 
    240.0303, 239.9912, 239.9521, 239.9521, 239.9131, 239.874,
  240.4603, 240.4212, 240.3822, 240.3431, 240.2649, 240.2258, 240.1867, 
    240.1476, 240.1085, 240.0694, 239.9912, 239.9521, 239.9131, 239.874, 
    239.8349, 239.7958, 239.7176, 239.6785, 239.6394, 239.6003,
  240.4603, 240.3822, 240.3431, 240.2649, 240.2258, 240.1867, 240.1085, 
    240.0694, 240.0303, 239.9521, 239.9131, 239.874, 239.8349, 239.7567, 
    239.7176, 239.6785, 239.6394, 239.6003, 239.5612, 239.483,
  240.3431, 240.304, 240.2649, 240.1867, 240.1476, 240.1085, 240.0694, 
    240.0303, 239.9912, 239.9521, 239.9131, 239.874, 239.8349, 239.7958, 
    239.7958, 239.7567, 239.7176, 239.6785, 239.6394, 239.6003,
  240.2649, 240.2258, 240.1867, 240.1476, 240.1085, 240.0694, 240.0303, 
    239.9912, 239.9912, 239.9521, 239.9521, 239.9131, 239.874, 239.874, 
    239.8349, 239.8349, 239.7958, 239.7958, 239.7567, 239.7567,
  240.2258, 240.1476, 240.1085, 240.0694, 240.0303, 239.9912, 239.9912, 
    239.9521, 239.9131, 239.874, 239.874, 239.8349, 239.8349, 239.7958, 
    239.7567, 239.7567, 239.7176, 239.6785, 239.6785, 239.6394,
  240.1476, 240.1085, 240.0694, 240.0303, 239.9912, 239.9521, 239.9521, 
    239.9131, 239.874, 239.874, 239.8349, 239.8349, 239.7958, 239.7567, 
    239.7567, 239.7176, 239.6785, 239.6394, 239.6003, 239.5612,
  240.1867, 240.1476, 240.1476, 240.1085, 240.1085, 240.1085, 240.0694, 
    240.0694, 240.0694, 240.0303, 240.0303, 239.9912, 239.9521, 239.9131, 
    239.874, 239.8349, 239.7958, 239.7176, 239.6785, 239.6003,
  240.4603, 240.4603, 240.4603, 240.4603, 240.4603, 240.4212, 240.4212, 
    240.4212, 240.3822, 240.3431, 240.3431, 240.2649, 240.2258, 240.1867, 
    240.1085, 240.0303, 239.9521, 239.874, 239.7958, 239.6785,
  240.6949, 240.6949, 240.6949, 240.6558, 240.6558, 240.6558, 240.6558, 
    240.6167, 240.5776, 240.5385, 240.4994, 240.4212, 240.3431, 240.2649, 
    240.1867, 240.0694, 239.9912, 239.874, 239.7176, 239.6003,
  240.6949, 240.6949, 240.6558, 240.6558, 240.6167, 240.6167, 240.5776, 
    240.5385, 240.4994, 240.4212, 240.3431, 240.2649, 240.1867, 240.1085, 
    239.9912, 239.8349, 239.7176, 239.5612, 239.4049, 239.2094,
  240.5776, 240.5385, 240.5385, 240.4994, 240.4603, 240.4212, 240.3822, 
    240.3431, 240.2649, 240.1867, 240.1085, 240.0303, 239.9131, 239.7958, 
    239.6394, 239.483, 239.3267, 239.1312, 238.9358, 238.7403,
  240.3431, 240.304, 240.2649, 240.2258, 240.1867, 240.1476, 240.1085, 
    240.0303, 239.9521, 239.874, 239.7958, 239.6785, 239.5612, 239.4049, 
    239.2485, 239.0921, 238.8967, 238.7012, 238.4667, 238.2321,
  240.0694, 240.0303, 239.9521, 239.9131, 239.874, 239.8349, 239.7958, 
    239.7176, 239.6394, 239.5221, 239.4049, 239.2876, 239.1312, 238.9358, 
    238.7403, 238.5449, 238.3494, 238.1149, 237.8803, 237.6458,
  239.9521, 239.874, 239.8349, 239.7958, 239.7958, 239.7567, 239.6785, 
    239.6394, 239.5221, 239.4049, 239.2876, 239.0921, 238.8967, 238.7012, 
    238.4667, 238.193, 237.9585, 237.6848, 237.4112, 237.1376,
  239.6785, 239.6394, 239.6003, 239.5612, 239.5221, 239.5221, 239.483, 
    239.444, 239.3658, 239.2485, 239.0921, 238.9358, 238.7012, 238.4667, 
    238.193, 237.8803, 237.6067, 237.2939, 236.9812, 236.6685,
  239.4049, 239.3267, 239.2876, 239.2094, 239.1703, 239.1312, 239.0921, 
    239.014, 238.9358, 238.7794, 238.623, 238.4276, 238.2321, 237.9585, 
    237.6848, 237.3721, 237.0985, 236.7858, 236.473, 236.1603,
  239.2876, 239.2485, 239.1703, 239.1312, 239.0531, 239.014, 238.9358, 
    238.8185, 238.7012, 238.5058, 238.3103, 238.0367, 237.7239, 237.4112, 
    237.0985, 236.7858, 236.473, 236.1603, 235.8475, 235.5739,
  226.2393, 226.2393, 226.2393, 226.2393, 226.2393, 226.2393, 226.2393, 
    226.2393, 226.2393, 226.2393, 226.2393, 226.2393, 226.2393, 226.2393, 
    226.2393, 226.2393, 226.2393, 226.2393, 226.2393, 226.2393,
  226.8552, 226.8552, 226.8552, 226.8552, 226.8552, 226.8552, 226.8552, 
    226.8552, 226.8552, 226.8552, 226.8552, 226.8552, 226.8552, 226.8552, 
    226.8552, 226.8552, 226.8552, 226.8552, 226.8552, 226.8552,
  226.9872, 226.9872, 226.9872, 226.9432, 226.9432, 226.9432, 226.9432, 
    226.8992, 226.8992, 226.8992, 226.8992, 226.8992, 226.8552, 226.8552, 
    226.8552, 226.8552, 226.8112, 226.8112, 226.8112, 226.8112,
  226.6792, 226.6353, 226.6353, 226.5913, 226.5473, 226.5473, 226.5033, 
    226.4593, 226.4153, 226.4153, 226.3713, 226.3713, 226.3273, 226.2833, 
    226.2833, 226.2393, 226.1953, 226.1953, 226.1514, 226.1074,
  226.1953, 226.1514, 226.0634, 226.0194, 225.9754, 225.9314, 225.8874, 
    225.8434, 225.7994, 225.7554, 225.7114, 225.6674, 225.6234, 225.5795, 
    225.5355, 225.4915, 225.4475, 225.4035, 225.3595, 225.3595,
  225.6234, 225.5795, 225.5355, 225.4915, 225.4475, 225.4035, 225.3595, 
    225.3155, 225.3155, 225.2715, 225.2715, 225.2275, 225.2275, 225.2275, 
    225.1835, 225.1835, 225.1835, 225.1395, 225.1395, 225.1395,
  225.5355, 225.4915, 225.4475, 225.4475, 225.4475, 225.4035, 225.4035, 
    225.4475, 225.4475, 225.4475, 225.4475, 225.4915, 225.4915, 225.5355, 
    225.5355, 225.5795, 225.5795, 225.6234, 225.6234, 225.6234,
  225.9314, 225.8874, 225.8874, 225.9314, 225.9314, 225.9754, 225.9754, 
    226.0194, 226.0634, 226.1074, 226.1953, 226.2393, 226.2833, 226.3273, 
    226.3713, 226.3713, 226.4153, 226.4593, 226.4593, 226.5033,
  226.2833, 226.2833, 226.3273, 226.3273, 226.4153, 226.4593, 226.5033, 
    226.5913, 226.6353, 226.7232, 226.7672, 226.8552, 226.8992, 226.9432, 
    226.9872, 227.0312, 227.0312, 227.0312, 227.0312, 227.0312,
  226.5473, 226.5913, 226.6353, 226.6792, 226.7672, 226.8552, 226.9432, 
    227.0312, 227.1192, 227.2072, 227.2951, 227.3831, 227.4711, 227.5151, 
    227.5591, 227.6031, 227.6031, 227.6031, 227.6031, 227.5591,
  227.1632, 227.2072, 227.2951, 227.3831, 227.4711, 227.6031, 227.6911, 
    227.823, 227.955, 228.043, 228.175, 228.263, 228.3069, 228.3949, 
    228.4389, 228.4389, 228.4389, 228.4389, 228.3949, 228.3509,
  227.867, 227.955, 228.087, 228.2189, 228.3509, 228.4829, 228.6589, 
    228.7908, 228.9228, 229.0108, 229.1428, 229.1868, 229.2747, 229.3187, 
    229.3187, 229.2747, 229.2747, 229.1868, 229.0988, 229.0108,
  228.5269, 228.6589, 228.7908, 228.9668, 229.1428, 229.2747, 229.4507, 
    229.5827, 229.7147, 229.8466, 229.9346, 229.9786, 229.9786, 229.9786, 
    229.9346, 229.8466, 229.7147, 229.5827, 229.4067, 229.2308,
  229.0108, 229.1428, 229.2747, 229.4507, 229.6267, 229.8027, 229.9786, 
    230.1546, 230.2866, 230.3745, 230.4625, 230.5065, 230.5065, 230.4185, 
    230.3306, 230.1986, 230.0226, 229.8027, 229.5827, 229.3187,
  229.2747, 229.3627, 229.4947, 229.6267, 229.8027, 229.9786, 230.1546, 
    230.3306, 230.4625, 230.5505, 230.5945, 230.6385, 230.5945, 230.5065, 
    230.3745, 230.1986, 230.0226, 229.7587, 229.4947, 229.2308,
  229.6267, 229.7587, 229.8906, 230.0226, 230.1546, 230.2866, 230.4185, 
    230.5505, 230.6385, 230.6825, 230.7265, 230.6825, 230.5945, 230.5065, 
    230.3306, 230.1106, 229.8906, 229.6707, 229.3627, 229.0988,
  230.0226, 230.1546, 230.3306, 230.5065, 230.6825, 230.8145, 230.9464, 
    231.0784, 231.1664, 231.1664, 231.1664, 231.0784, 230.9025, 230.7265, 
    230.5065, 230.2426, 229.9346, 229.6707, 229.3627, 229.0548,
  230.2866, 230.4185, 230.5945, 230.7705, 230.9904, 231.1664, 231.2984, 
    231.4303, 231.5183, 231.5183, 231.4743, 231.3864, 231.2104, 230.9904, 
    230.7265, 230.4625, 230.1546, 229.8027, 229.4947, 229.1428,
  230.8585, 230.9904, 231.1224, 231.2984, 231.4743, 231.5623, 231.6503, 
    231.7383, 231.7383, 231.7383, 231.6943, 231.5623, 231.3864, 231.1664, 
    230.9025, 230.5945, 230.3306, 230.0226, 229.7147, 229.4067,
  231.9142, 232.0462, 232.1782, 232.3542, 232.4422, 232.5301, 232.5741, 
    232.5741, 232.5301, 232.3982, 232.2222, 231.9582, 231.6503, 231.3424, 
    231.0344, 230.7705, 230.4625, 230.1546, 229.8466, 229.5387,
  218.8314, 218.8314, 218.8314, 218.8314, 218.8314, 218.8314, 218.8314, 
    218.8314, 218.8314, 218.8314, 218.8314, 218.8314, 218.8314, 218.8314, 
    218.8799, 218.8799, 218.8799, 218.8799, 218.8799, 218.8799,
  219.1225, 219.171, 219.171, 219.171, 219.171, 219.171, 219.171, 219.171, 
    219.171, 219.2195, 219.2195, 219.2195, 219.2195, 219.2195, 219.2195, 
    219.2195, 219.2195, 219.2195, 219.2195, 219.2195,
  218.9769, 218.9769, 218.9769, 218.9769, 218.9769, 218.9769, 218.9769, 
    218.9284, 218.9284, 218.9284, 218.9284, 218.9284, 218.9284, 218.9284, 
    218.9284, 218.9284, 218.9284, 218.9284, 218.9284, 218.9284,
  218.7829, 218.7829, 218.7344, 218.6859, 218.6373, 218.6373, 218.5888, 
    218.5403, 218.5403, 218.4918, 218.4433, 218.4433, 218.3948, 218.3463, 
    218.3463, 218.2977, 218.2492, 218.2492, 218.2007, 218.1522,
  218.6373, 218.5403, 218.4433, 218.3948, 218.2977, 218.2492, 218.1522, 
    218.1037, 218.0552, 217.9582, 217.9096, 217.8611, 217.8126, 217.7156, 
    217.6671, 217.6186, 217.5701, 217.5215, 217.473, 217.4245,
  218.0552, 217.9582, 217.8611, 217.7641, 217.6671, 217.6186, 217.5701, 
    217.473, 217.4245, 217.376, 217.3275, 217.279, 217.279, 217.2305, 
    217.1819, 217.1819, 217.1334, 217.1334, 217.0849, 217.0364,
  218.0067, 217.9096, 217.8126, 217.7641, 217.7156, 217.6671, 217.6671, 
    217.6186, 217.6186, 217.6186, 217.6186, 217.6186, 217.6186, 217.6186, 
    217.6186, 217.6671, 217.6671, 217.7156, 217.7156, 217.7641,
  218.6373, 218.5403, 218.4918, 218.4433, 218.4433, 218.3948, 218.3948, 
    218.3948, 218.4433, 218.4918, 218.4918, 218.5403, 218.5888, 218.6373, 
    218.6859, 218.7344, 218.7829, 218.8314, 218.8799, 218.9284,
  218.6373, 218.5888, 218.5403, 218.5403, 218.5403, 218.5888, 218.5888, 
    218.6373, 218.6859, 218.7344, 218.8314, 218.8799, 218.9284, 219.0255, 
    219.074, 219.1225, 219.2195, 219.268, 219.268, 219.3165,
  218.4918, 218.4433, 218.4433, 218.4433, 218.4918, 218.5403, 218.6373, 
    218.6859, 218.7829, 218.8799, 218.9769, 219.1225, 219.2195, 219.3165, 
    219.365, 219.4621, 219.5106, 219.5591, 219.6076, 219.6076,
  218.8799, 218.8314, 218.8799, 218.9284, 219.0255, 219.1225, 219.2195, 
    219.3165, 219.4621, 219.6076, 219.7046, 219.8502, 219.9472, 220.0442, 
    220.1413, 220.2383, 220.2868, 220.2868, 220.2868, 220.2868,
  219.4136, 219.4621, 219.5591, 219.6561, 219.8017, 219.9472, 220.0927, 
    220.2383, 220.4323, 220.5779, 220.6749, 220.8204, 220.9175, 220.966, 
    221.0145, 221.0145, 221.0145, 220.966, 220.9175, 220.8204,
  219.8987, 219.9957, 220.1413, 220.3353, 220.5294, 220.7234, 220.9175, 
    221.1115, 221.3056, 221.4511, 221.5966, 221.6937, 221.7422, 221.7907, 
    221.7422, 221.6937, 221.5966, 221.4511, 221.3056, 221.1115,
  220.4809, 220.6264, 220.7719, 220.966, 221.16, 221.4026, 221.6452, 
    221.8392, 222.0333, 222.2273, 222.3729, 222.4699, 222.5184, 222.4699, 
    222.4214, 222.3244, 222.1788, 221.9362, 221.7422, 221.4511,
  220.7719, 220.9175, 221.063, 221.3056, 221.4996, 221.7422, 221.9848, 
    222.2273, 222.4214, 222.6154, 222.761, 222.858, 222.9065, 222.858, 
    222.8095, 222.664, 222.5184, 222.2758, 222.0333, 221.7422,
  221.0145, 221.16, 221.3541, 221.5966, 221.8392, 222.0818, 222.3244, 
    222.5669, 222.761, 222.9065, 223.0521, 223.1006, 223.1006, 223.0521, 
    222.9065, 222.761, 222.5184, 222.2758, 221.9848, 221.6452,
  221.4996, 221.6452, 221.8877, 222.1788, 222.4699, 222.761, 223.0035, 
    223.1976, 223.3916, 223.4887, 223.5372, 223.4887, 223.3916, 223.2461, 
    223.0035, 222.761, 222.4214, 222.1303, 221.7907, 221.4026,
  221.5481, 221.7422, 221.9848, 222.2758, 222.5669, 222.9065, 223.1491, 
    223.3916, 223.5372, 223.6342, 223.6827, 223.5857, 223.4402, 223.2461, 
    223.0035, 222.7125, 222.3729, 222.0333, 221.6452, 221.3056,
  221.5966, 221.8392, 222.1303, 222.4214, 222.7125, 222.955, 223.1976, 
    223.3431, 223.4402, 223.4887, 223.4887, 223.3916, 223.2461, 223.0521, 
    222.8095, 222.5184, 222.1788, 221.8392, 221.4511, 221.1115,
  222.5669, 222.761, 223.0035, 223.1976, 223.3431, 223.5372, 223.6827, 
    223.7798, 223.8283, 223.7798, 223.6827, 223.4887, 223.2461, 222.955, 
    222.664, 222.3244, 221.9362, 221.5481, 221.1115, 220.7234 ;
}
