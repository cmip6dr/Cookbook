netcdf hurs_Amon_exAA05_decadal1981_r1i1p1_198201-199112_box {
dimensions:
	lon = 20 ;
	bnds = 2 ;
	lat = 20 ;
	time = UNLIMITED ; // (4 currently)
variables:
	double lon(lon) ;
		lon:standard_name = "longitude" ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:axis = "X" ;
		lon:bounds = "lon_bnds" ;
	double lon_bnds(lon, bnds) ;
	double lat(lat) ;
		lat:standard_name = "latitude" ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:axis = "Y" ;
		lat:bounds = "lat_bnds" ;
	double lat_bnds(lat, bnds) ;
	double height ;
		height:standard_name = "height" ;
		height:long_name = "height" ;
		height:units = "m" ;
		height:positive = "up" ;
		height:axis = "Z" ;
	double time(time) ;
		time:standard_name = "time" ;
		time:long_name = "time" ;
		time:bounds = "time_bnds" ;
		time:units = "days since 1982-1-1 00:00:00" ;
		time:calendar = "365_day" ;
		time:axis = "T" ;
	double time_bnds(time, bnds) ;
	float hurs(time, lat, lon) ;
		hurs:standard_name = "relative_humidity" ;
		hurs:long_name = "Near-Surface Relative Humidity" ;
		hurs:units = "%" ;
		hurs:grid_type = "gaussian" ;
		hurs:coordinates = "height" ;
		hurs:_FillValue = 1.e+20f ;
		hurs:missing_value = 1.e+20f ;
		hurs:comment = "This is the relative humidity with respect to liquid water for T> 0 C, and with respect to ice for T<0 C." ;
		hurs:original_name = "HURS" ;
		hurs:cell_methods = "time: mean (interval: 20 mintues)" ;
		hurs:history = "2012-08-15T07:31:53Z altered by CMOR: Treated scalar dimension: \'height\'." ;
		hurs:associated_files = "baseURL: http://cmip-pcmdi.llnl.gov/CMIP5/dataLocation gridspecFile: gridspec_atmos_fx_bcc-csm1-1_decadal1981_r0i0p0.nc areacella: areacella_fx_bcc-csm1-1_decadal1981_r0i0p0.nc" ;

// global attributes:
		:CDI = "Climate Data Interface version ?? (http://mpimet.mpg.de/cdi)" ;
		:Conventions = "CF-1.4" ;
		:history = "reset by cdo to create anonymous sample file" ;
		:source = "201707_compliance_checker_evaluation/work/p1.py" ;
		:institution = "CEDA" ;
		:institute_id = "CEDA" ;
		:experiment_id = "decadal1981" ;
		:model_id = "exAA05" ;
		:forcing = "Nat Ant GHG SD Oz Sl Vl SS Ds BC OC" ;
		:parent_experiment_id = "historical" ;
		:parent_experiment_rip = "r1i1p1" ;
		:branch_time = 1981. ;
		:contact = "none" ;
		:comment = "this is a sample file with known metadata errors" ;
		:initialization_method = 1 ;
		:physics_version = 1 ;
		:tracking_id = "37994f26-9f35-4e36-b539-8c9cdfa36487" ;
		:product = "output" ;
		:experiment = "10- or 30-year run initialized in year 1981" ;
		:frequency = "mon" ;
		:creation_date = "2012-08-15T07:31:54Z" ;
		:project_id = "CMIP5" ;
		:table_id = "Table Amon (11 April 2011) 1cfdc7322cf2f4a32614826fab42c1ab" ;
		:title = "Dummy file with known metadata errors" ;
		:parent_experiment = "historical" ;
		:modeling_realm = "atmos" ;
		:realization = 1 ;
		:cmor_version = "2.5.6" ;
		:CDO = "Climate Data Operators version 1.7.0 (http://mpimet.mpg.de/cdo)" ;
data:

 lon = 0, 2.8125, 5.625, 8.4375, 11.25, 14.0625, 16.875, 19.6875, 22.5, 
    25.3125, 28.125, 30.9375, 33.75, 36.5625, 39.375, 42.1875, 45, 47.8125, 
    50.625, 53.4375 ;

 lon_bnds =
  -1.40625, 1.40625,
  1.40625, 4.21875,
  4.21875, 7.03125,
  7.03125, 9.84375,
  9.84375, 12.65625,
  12.65625, 15.46875,
  15.46875, 18.28125,
  18.28125, 21.09375,
  21.09375, 23.90625,
  23.90625, 26.71875,
  26.71875, 29.53125,
  29.53125, 32.34375,
  32.34375, 35.15625,
  35.15625, 37.96875,
  37.96875, 40.78125,
  40.78125, 43.59375,
  43.59375, 46.40625,
  46.40625, 49.21875,
  49.21875, 52.03125,
  52.03125, 54.84375 ;

 lat = -87.8637988392326, -85.0965269883174, -82.3129129478863, 
    -79.5256065726594, -76.7368996803683, -73.9475151539897, 
    -71.1577520115873, -68.3677561083132, -65.5776070108278, 
    -62.7873517989631, -59.9970201084913, -57.2066315276432, 
    -54.4161995260862, -51.6257336749383, -48.8352409662506, 
    -46.0447266311017, -43.2541946653509, -40.463648178115, 
    -37.6730896290453, -34.8825209937735 ;

 lat_bnds =
  -87.8637988392326, -86.480162913775,
  -86.480162913775, -83.7047199681018,
  -83.7047199681018, -80.9192597602729,
  -80.9192597602729, -78.1312531265139,
  -78.1312531265139, -75.342207417179,
  -75.342207417179, -72.5526335827885,
  -72.5526335827885, -69.7627540599503,
  -69.7627540599503, -66.9726815595705,
  -66.9726815595705, -64.1824794048954,
  -64.1824794048954, -61.3921859537272,
  -61.3921859537272, -58.6018258180673,
  -58.6018258180673, -55.8114155268647,
  -55.8114155268647, -53.0209666005122,
  -53.0209666005122, -50.2304873205944,
  -50.2304873205944, -47.4399837986761,
  -47.4399837986761, -44.6494606482263,
  -44.6494606482263, -41.858921421733,
  -41.858921421733, -39.0683689035802,
  -39.0683689035802, -36.2778053114094,
  -36.2778053114094, -33.4872324377587 ;

 height = 2 ;

 time = 15.5, 45, 74.5, 105 ;

 time_bnds =
  0, 31,
  31, 59,
  59, 90,
  90, 120 ;

 hurs =
  93.4809, 93.74128, 93.9556, 94.03909, 94.47622, 94.65362, 94.82246, 
    95.1601, 93.7446, 94.10422, 94.16572, 94.11856, 94.13337, 94.49639, 
    94.70043, 94.81069, 93.98279, 94.30159, 94.16895, 94.13051,
  88.7273, 89.54988, 90.32349, 91.12242, 92.00128, 92.69608, 93.63831, 
    94.38155, 91.08723, 91.9362, 92.52862, 93.34216, 93.92194, 94.5956, 
    94.90078, 95.31381, 93.43739, 94.07809, 94.69255, 95.03079,
  83.48702, 84.99387, 86.29594, 87.70504, 88.8302, 89.77134, 91.012, 
    92.43107, 88.70104, 89.85878, 90.94014, 92.18761, 92.81371, 93.41303, 
    93.52509, 94.11451, 92.28455, 92.71619, 93.31631, 93.52835,
  84.69096, 86.19128, 87.67854, 89.19056, 90.50443, 91.71695, 92.53498, 
    93.33336, 90.69014, 91.27824, 91.97832, 92.61449, 93.1025, 93.40945, 
    93.54196, 93.37686, 93.75618, 93.67755, 93.39366, 93.51973,
  83.67885, 86.10898, 88.38322, 90.29052, 91.65009, 92.62195, 93.09725, 
    93.88835, 91.5418, 91.3267, 91.20734, 91.85376, 92.48512, 92.65701, 
    92.91588, 92.77927, 96.84536, 96.78885, 96.07845, 95.499,
  82.51562, 84.88831, 86.97651, 88.77648, 89.76414, 90.14468, 90.25821, 
    90.01252, 85.492, 85.72311, 86.30702, 87.01633, 88.00871, 89.5621, 
    91.02483, 92.61087, 98.50533, 98.64861, 98.5509, 98.17497,
  89.68507, 86.78841, 86.6087, 86.84266, 86.71143, 86.51164, 86.33993, 
    85.93306, 77.86455, 77.40113, 77.35551, 79.10056, 81.01414, 85.01857, 
    84.12335, 87.63353, 94.95633, 96.56116, 97.33598, 97.23394,
  93.43623, 92.90776, 91.67722, 90.48186, 89.21488, 88.15541, 87.04222, 
    85.63926, 77.28253, 75.64349, 75.49283, 78.94083, 78.86671, 79.91819, 
    70.37437, 74.3143, 78.09537, 93.66832, 94.12508, 95.66349,
  87.42145, 88.93051, 90.46446, 91.42157, 91.6532, 91.33952, 90.35046, 
    88.95781, 84.75066, 83.16238, 82.43893, 82.44582, 83.63319, 84.69102, 
    85.57793, 86.90664, 88.29635, 88.45477, 91.93355, 94.33942,
  84.33488, 86.3585, 88.88643, 91.39141, 92.21031, 91.9331, 91.31547, 
    90.97707, 90.83997, 90.39748, 90.02382, 89.0844, 88.53478, 88.39187, 
    88.94681, 89.19878, 89.81826, 91.08138, 92.13571, 92.45863,
  81.94168, 82.978, 84.72486, 87.94966, 90.65647, 91.54073, 91.38587, 
    91.50724, 92.07696, 92.36807, 92.84383, 92.41033, 91.17633, 90.46159, 
    90.12606, 89.69244, 89.76153, 89.78741, 90.41199, 91.27546,
  82.42509, 82.66344, 83.24526, 85.00698, 86.61463, 86.95371, 86.59507, 
    87.69249, 90.12206, 91.88249, 92.80717, 92.99869, 92.13709, 91.56483, 
    91.09361, 89.98956, 89.55358, 89.58495, 89.884, 90.68936,
  85.83164, 85.98697, 86.30321, 86.7794, 86.6998, 84.66866, 81.7151, 
    81.01419, 83.48742, 86.76139, 89.18749, 90.869, 91.45655, 91.09351, 
    91.39294, 91.30672, 90.09115, 88.65224, 88.784, 89.37923,
  82.37218, 83.16448, 83.78975, 84.20922, 83.2514, 81.95366, 81.78837, 
    82.77064, 84.525, 86.61893, 87.79867, 88.67591, 89.51363, 90.13094, 
    91.13078, 91.47941, 89.81043, 88.1453, 87.87795, 89.09147,
  75.86752, 75.09309, 75.2433, 75.39053, 75.22278, 76.72486, 80.25311, 
    83.74046, 86.40416, 87.6395, 88.04431, 88.57058, 89.66587, 90.52764, 
    90.9056, 91.11395, 90.21503, 89.09438, 89.44652, 90.82539,
  73.35105, 72.47985, 72.89262, 74.36884, 76.2441, 78.83097, 82.01714, 
    84.33385, 86.53508, 88.42753, 89.38844, 89.757, 90.1792, 90.89043, 
    91.0164, 90.70487, 89.87632, 89.47755, 90.27154, 90.51128,
  76.63313, 77.2861, 78.97208, 80.56419, 81.63042, 82.18461, 82.20987, 
    82.44176, 84.14093, 86.33018, 88.35344, 89.31207, 89.28953, 89.42931, 
    89.32444, 88.2574, 86.47741, 85.4045, 84.93102, 84.50637,
  83.00284, 82.76088, 82.8689, 81.82735, 80.72785, 79.71549, 79.37939, 
    78.76436, 74.75816, 73.10941, 74.78475, 78.0412, 80.88372, 82.72076, 
    84.10639, 84.26265, 82.52142, 79.37403, 77.83792, 78.10139,
  81.83013, 80.74139, 79.26865, 77.1935, 75.92776, 76.23385, 75.38225, 
    69.07002, 63.52311, 61.11913, 61.72075, 65.10432, 69.99793, 74.59365, 
    78.36984, 79.33351, 78.0505, 77.30078, 78.44856, 80.42095,
  73.47881, 72.02462, 70.44322, 69.69109, 69.98117, 70.39768, 67.90502, 
    63.09711, 60.43573, 58.8373, 59.27411, 63.01844, 70.89108, 76.50346, 
    78.50382, 78.2642, 78.4737, 79.86833, 81.52776, 82.52912,
  91.05083, 91.30476, 91.53485, 92.02209, 92.18385, 92.56113, 92.62751, 
    93.08926, 91.88125, 92.40703, 92.5981, 92.64035, 92.99768, 92.64845, 
    93.51599, 93.89808, 92.04053, 93.13046, 92.65516, 93.22881,
  86.96413, 87.80626, 88.72099, 89.57648, 90.3923, 91.21534, 92.04106, 
    92.90271, 89.44534, 90.34664, 91.18976, 92.07103, 92.96951, 93.7209, 
    94.42259, 95.10692, 93.32484, 94.06727, 94.6227, 94.98904,
  85.80513, 87.10407, 88.54015, 89.99532, 91.11778, 92.29962, 93.42702, 
    94.41877, 90.26347, 91.3447, 92.29098, 93.48471, 94.67207, 95.65806, 
    96.47842, 97.24012, 95.63651, 96.28072, 96.89655, 97.20786,
  85.95926, 87.22572, 88.69738, 90.30405, 91.83503, 92.93233, 94.13572, 
    95.26557, 93.02795, 94.30644, 95.31511, 95.90936, 96.54295, 97.02541, 
    97.50476, 97.7431, 98.66412, 98.55714, 98.53976, 97.77951,
  84.73331, 86.33834, 88.74374, 90.77811, 92.45103, 93.38811, 94.29533, 
    95.24791, 94.00957, 94.55647, 94.90408, 95.08174, 95.35646, 96.20399, 
    96.47029, 96.29651, 99.09619, 98.84468, 98.37006, 97.46123,
  84.39301, 86.8561, 88.84941, 90.42979, 91.79298, 92.48118, 92.73416, 
    92.78191, 88.05251, 88.12733, 88.48933, 88.75777, 89.77502, 90.84673, 
    91.97835, 93.42875, 98.78717, 98.84388, 98.49764, 98.00574,
  88.28484, 85.12112, 84.33315, 84.39015, 84.37801, 84.40788, 84.34162, 
    84.17943, 76.47164, 75.87708, 75.25665, 74.02428, 76.02343, 84.70475, 
    85.37189, 84.09641, 92.42211, 95.36664, 96.6904, 97.2202,
  70.56541, 68.4983, 67.41721, 66.8833, 67.7931, 69.21661, 69.8529, 69.42115, 
    63.17681, 62.5233, 62.89027, 67.26984, 66.06211, 65.23525, 55.66279, 
    58.71144, 67.86268, 87.54339, 86.85458, 88.93345,
  68.84487, 68.51212, 69.35588, 71.91167, 74.11705, 75.94108, 76.46138, 
    75.37688, 71.65511, 70.68373, 70.22173, 70.43938, 71.64607, 72.97045, 
    74.19555, 75.15436, 74.11209, 71.4112, 75.65611, 78.24518,
  76.204, 75.76051, 76.30462, 78.38274, 80.0094, 80.87751, 81.61044, 
    81.53532, 81.66994, 81.50655, 81.2676, 81.04417, 81.54856, 82.12254, 
    81.42691, 81.53082, 82.43788, 82.96621, 83.54175, 83.96078,
  80.23288, 79.93113, 79.55199, 80.25504, 81.74779, 82.56519, 82.99827, 
    83.67518, 84.84621, 85.20068, 86.04611, 86.85261, 87.18818, 86.70637, 
    85.09091, 83.79376, 83.47128, 83.66501, 84.92827, 87.11862,
  80.3205, 80.81688, 80.38798, 80.2877, 80.36696, 80.49259, 80.68171, 
    81.90107, 84.04259, 86.0901, 87.90427, 89.13175, 89.38041, 88.99027, 
    87.82668, 86.39554, 85.45226, 85.01891, 85.1569, 85.85855,
  82.61204, 84.35664, 84.58595, 83.7952, 83.19865, 82.12931, 80.47408, 
    80.31496, 81.63389, 84.10897, 86.23838, 88.20938, 89.64275, 90.14081, 
    90.22598, 89.43638, 87.71576, 85.99191, 85.64497, 86.32988,
  77.52943, 80.00568, 81.99464, 82.82799, 82.7672, 81.90527, 81.63331, 
    82.93295, 84.85116, 86.85659, 88.73515, 90.06676, 91.00152, 91.6852, 
    92.33061, 92.27951, 91.1763, 90.12089, 90.0131, 90.05972,
  70.85555, 71.13307, 72.69428, 75.08057, 76.58379, 77.37475, 79.43566, 
    82.78063, 85.86054, 88.28426, 90.07277, 91.17024, 91.87083, 91.45269, 
    90.72025, 90.61872, 90.62669, 90.56753, 90.9033, 91.29102,
  67.00684, 67.09906, 68.57079, 71.75898, 74.98229, 77.92363, 81.4397, 
    83.80692, 85.61021, 87.91116, 89.82823, 90.51535, 90.31052, 89.72369, 
    89.45454, 89.80968, 89.86005, 89.7135, 90.07793, 89.7205,
  67.42973, 69.64367, 73.03672, 76.33788, 78.47476, 80.10015, 81.0109, 
    81.44915, 82.62988, 84.73471, 86.24037, 86.77477, 86.97071, 87.5002, 
    87.86768, 87.51228, 86.24092, 84.8092, 83.44328, 81.98793,
  71.84314, 73.90975, 76.41698, 77.60235, 77.50567, 77.15674, 76.7172, 
    76.34422, 73.36298, 72.05531, 73.5601, 76.21287, 79.43002, 81.82706, 
    82.31962, 81.0184, 78.15611, 74.86246, 73.23536, 72.86601,
  72.87029, 73.06731, 73.01364, 72.42223, 71.79234, 72.95309, 72.38346, 
    67.12737, 64.14597, 63.28709, 64.52564, 67.76785, 72.1254, 74.02386, 
    73.94988, 72.74982, 70.37342, 69.23614, 70.56975, 72.32249,
  66.57248, 65.85196, 64.97097, 64.76868, 66.37942, 68.13031, 66.52633, 
    63.15863, 64.16334, 65.31944, 65.01894, 65.8837, 69.25704, 71.14582, 
    70.45712, 69.66892, 70.43227, 72.44795, 74.49334, 76.20102,
  92.22964, 92.43774, 92.63062, 92.8927, 93.19102, 93.51788, 93.97072, 
    94.11161, 92.57564, 92.95654, 92.68084, 92.93453, 92.90622, 93.64265, 
    93.20396, 93.64107, 92.85706, 93.42496, 93.58959, 94.07526,
  86.53026, 87.48244, 88.50666, 89.69047, 90.90907, 91.94442, 92.98344, 
    94.28337, 91.34309, 92.40143, 93.23909, 93.97713, 94.6262, 95.10246, 
    95.59241, 96.23475, 94.76723, 95.52543, 96.14085, 96.77498,
  86.57798, 88.27718, 90.18165, 92.02053, 93.36674, 94.7112, 95.64027, 
    96.24773, 92.06914, 93.2021, 94.23994, 95.49935, 96.77421, 97.63377, 
    97.98104, 98.39999, 97.01608, 97.34422, 97.65852, 98.02956,
  85.57472, 87.42229, 89.42072, 91.31242, 92.87572, 94.0182, 94.81004, 
    95.25046, 92.9412, 93.63285, 94.24619, 94.66399, 95.5916, 96.98648, 
    97.69051, 97.93504, 98.9244, 99.30836, 99.28754, 99.01913,
  79.8897, 81.06566, 83.05697, 84.85406, 86.71394, 88.3033, 89.21417, 
    90.49871, 89.98582, 90.96175, 90.5547, 91.20617, 91.58131, 92.33372, 
    92.52147, 92.46666, 95.38915, 95.59892, 95.88333, 95.71642,
  81.32919, 83.57585, 85.60041, 87.10515, 87.96142, 88.2849, 88.83413, 
    89.01068, 84.51334, 84.6098, 85.05444, 85.95848, 86.76998, 87.46896, 
    87.9019, 88.61512, 94.58236, 95.06998, 95.14769, 94.7646,
  88.07307, 86.59868, 86.58923, 85.98232, 87.31383, 89.03308, 87.69571, 
    86.28378, 78.07515, 77.42992, 76.50029, 75.31867, 77.60992, 84.57999, 
    88.4496, 83.90228, 90.68993, 92.63293, 93.92556, 94.3019,
  66.82751, 64.60086, 62.82958, 61.60794, 63.41624, 65.40393, 63.58063, 
    61.02935, 54.88851, 52.43182, 52.38718, 59.72296, 63.81407, 71.09298, 
    73.98959, 77.97992, 85.19641, 87.71232, 85.54469, 85.85326,
  73.13551, 71.02815, 69.26849, 68.40961, 68.70718, 70.467, 72.87477, 
    74.51218, 72.79417, 72.56232, 72.75586, 73.20984, 73.98312, 74.24403, 
    72.93912, 70.91954, 68.17037, 66.61717, 71.47506, 76.72422,
  79.34602, 78.66451, 78.3548, 77.70069, 76.63519, 76.07726, 76.30894, 
    76.85977, 77.66917, 78.23744, 78.81143, 79.5592, 80.23734, 80.9165, 
    81.75278, 81.83458, 81.53395, 81.31597, 81.78459, 81.8632,
  82.1837, 81.05145, 80.16758, 79.96313, 79.35477, 78.85178, 79.16402, 
    79.59003, 80.19248, 80.37486, 80.93359, 81.53082, 82.25062, 83.12988, 
    83.54334, 83.05065, 82.54458, 82.45341, 83.38203, 85.05447,
  82.27977, 81.84331, 81.39489, 81.61255, 81.11818, 80.31812, 79.75488, 
    80.21078, 81.15015, 82.00865, 82.57651, 82.95551, 83.45312, 84.68269, 
    85.90909, 85.93105, 85.15443, 84.02096, 83.69626, 84.02985,
  83.19819, 84.77756, 85.29516, 85.23341, 84.3204, 81.84599, 78.9753, 
    78.56066, 80.26664, 82.85178, 84.57373, 85.59086, 86.2681, 87.16847, 
    88.62134, 89.42458, 88.9723, 87.42092, 86.10884, 85.40966,
  77.55661, 78.20733, 78.97232, 78.85659, 77.29427, 75.32452, 73.60342, 
    73.67761, 76.62664, 80.55087, 83.18075, 85.25797, 87.23463, 89.3175, 
    91.49753, 91.87869, 91.04417, 90.20111, 89.73278, 89.18158,
  72.69135, 71.18095, 70.91507, 71.17534, 70.98412, 71.0764, 71.73852, 
    74.35057, 78.77151, 82.15887, 84.43987, 86.56584, 88.47732, 90.17076, 
    91.45909, 91.71172, 91.01821, 90.18664, 90.21486, 90.02959,
  71.88069, 70.26759, 69.84135, 70.97539, 72.88988, 75.61446, 78.73995, 
    81.53966, 83.13571, 84.78057, 86.86706, 88.44273, 89.37089, 89.90425, 
    89.52814, 88.78856, 87.91721, 86.92907, 87.05277, 86.4493,
  75.1648, 75.33139, 76.83544, 78.9208, 80.75966, 81.75249, 81.45548, 
    80.67786, 81.05466, 83.27165, 85.56857, 86.81513, 87.19731, 87.20964, 
    85.99469, 84.66291, 83.5312, 82.70512, 82.69513, 82.53698,
  80.13885, 80.93002, 82.51959, 82.78947, 81.56464, 79.74812, 78.35667, 
    76.45396, 71.82506, 70.24403, 72.7714, 76.51721, 79.09177, 80.22096, 
    81.24654, 81.64393, 80.49542, 79.13195, 78.72643, 78.86671,
  78.32669, 78.63792, 78.58054, 76.83755, 75.471, 75.81986, 74.33036, 
    67.22467, 61.09481, 59.61237, 61.09739, 64.24065, 68.30055, 72.31342, 
    76.53555, 78.25968, 77.88239, 77.30264, 77.3987, 77.07419,
  68.94539, 68.68242, 67.90125, 67.52906, 68.38454, 68.82463, 66.44341, 
    64.24481, 64.48137, 66.51134, 66.76366, 67.10056, 71.16967, 76.8642, 
    79.77894, 78.94858, 78.6658, 79.55561, 79.34438, 78.17169,
  92.54141, 93.03654, 93.52762, 93.84403, 94.29354, 94.51123, 94.85713, 
    95.37252, 93.90202, 94.31615, 94.88012, 95.2742, 95.43367, 95.5916, 
    95.6601, 95.76815, 94.76352, 94.81911, 95.11162, 94.88686,
  88.01664, 89.33185, 90.5452, 91.72334, 93.03945, 94.02189, 94.6624, 
    95.15916, 91.48368, 92.13939, 92.6049, 93.2338, 94.24551, 95.44672, 
    96.71396, 97.30254, 96.08929, 97.30815, 98.098, 98.56557,
  90.94303, 92.52785, 93.59134, 94.15833, 94.02104, 94.04562, 94.29615, 
    95.22523, 92.14843, 93.13724, 94.34363, 95.3501, 95.84255, 96.49215, 
    97.14639, 97.7093, 96.85003, 96.86707, 98.12727, 98.75555,
  88.27318, 90.09724, 90.99214, 92.27362, 93.60272, 94.15263, 94.1814, 
    93.75691, 92.58743, 94.21455, 95.44579, 95.48254, 97.53008, 98.88947, 
    99.46278, 99.73093, 99.77509, 99.8382, 99.89862, 99.71155,
  87.89031, 90.40994, 91.82758, 92.53615, 90.4079, 89.04392, 86.26049, 
    84.59306, 84.01423, 84.81204, 87.06075, 90.74068, 92.94947, 94.75008, 
    96.19665, 97.18544, 98.77139, 98.6069, 98.57997, 98.00607,
  83.8903, 84.92136, 85.39373, 85.37511, 84.69858, 83.02608, 82.80133, 
    82.95575, 79.49889, 80.70763, 82.39478, 84.50827, 86.53953, 88.32211, 
    89.75426, 90.74025, 97.06171, 97.45334, 97.07273, 96.55278,
  90.88854, 89.76771, 89.11231, 88.62409, 87.96299, 88.64448, 89.22742, 
    89.59662, 83.00499, 84.28205, 85.38667, 75.99948, 78.06296, 86.1804, 
    91.22605, 85.66981, 91.63414, 93.50183, 94.56201, 95.41918,
  68.94415, 66.33955, 64.29183, 65.86238, 68.57698, 72.97327, 75.46369, 
    75.94781, 70.16953, 71.42984, 75.55386, 78.06153, 82.2213, 89.04475, 
    92.60138, 93.229, 94.92187, 93.98281, 90.93874, 89.7681,
  71.95364, 69.37602, 67.37003, 65.48115, 64.44978, 64.15454, 64.02914, 
    64.00714, 62.10726, 62.3767, 63.09856, 64.20993, 65.98297, 68.32056, 
    69.56511, 70.84837, 74.83064, 81.55328, 86.19711, 88.44236,
  80.79776, 81.13727, 80.99896, 80.06807, 78.51117, 76.4956, 74.8095, 
    73.18134, 72.48692, 72.22964, 72.51437, 73.08861, 73.94782, 75.33536, 
    76.24101, 76.79229, 77.74096, 77.86268, 77.6832, 76.9064,
  82.41901, 82.753, 82.95709, 83.02888, 82.5001, 81.62798, 80.52926, 
    79.42319, 79.03169, 78.65395, 78.60709, 78.77505, 79.4987, 80.38777, 
    80.64737, 80.33028, 80.24097, 79.32241, 78.44655, 78.81319,
  82.85352, 83.37037, 83.26756, 83.29868, 82.87095, 81.83881, 81.79357, 
    83.27275, 85.26991, 85.91756, 85.69547, 85.26593, 85.25497, 85.41699, 
    85.35724, 84.64681, 83.86331, 82.14967, 80.87762, 80.50623,
  83.38592, 85.35951, 86.53141, 86.30074, 85.66002, 84.33922, 81.94282, 
    80.93518, 81.83748, 83.32011, 84.69791, 86.03635, 87.139, 87.7773, 
    88.77158, 89.18918, 88.49197, 86.56252, 84.66927, 82.93718,
  75.79934, 76.75446, 77.52898, 77.5277, 76.99945, 76.20707, 75.2501, 
    74.26753, 74.8577, 77.57658, 80.82764, 84.20567, 87.21058, 89.12047, 
    90.78375, 91.23209, 90.35426, 89.3278, 88.5433, 86.92542,
  69.21698, 68.35692, 68.80516, 69.58924, 70.05959, 70.75885, 71.75528, 
    73.23194, 77.27584, 82.16837, 86.12025, 88.95671, 90.60925, 90.88049, 
    90.78745, 90.44984, 89.46867, 88.44221, 88.83672, 89.24079,
  68.50562, 68.10552, 68.59997, 70.33549, 72.60332, 75.29845, 78.04709, 
    80.88697, 83.91629, 86.45277, 88.43858, 89.40572, 89.91223, 90.19718, 
    90.01281, 89.71179, 89.20315, 88.67767, 89.69603, 89.97243,
  71.52088, 73.22936, 75.69386, 78.65891, 81.17647, 82.8969, 83.16904, 
    82.24049, 81.93842, 83.45264, 86.2891, 87.97657, 88.5819, 88.9337, 
    88.85368, 88.32925, 87.61467, 86.53557, 86.01635, 85.59343,
  75.79662, 78.00786, 80.5469, 81.59884, 80.70174, 78.97758, 77.41759, 
    74.14724, 69.33091, 69.06882, 72.36685, 76.35325, 79.35719, 81.87857, 
    83.53662, 83.43586, 81.40395, 78.64791, 77.64761, 78.19087,
  75.40871, 75.86194, 75.55762, 73.83998, 72.1325, 71.50379, 69.34479, 
    62.2871, 58.01443, 56.88947, 57.08403, 58.79262, 62.98716, 68.70476, 
    73.22769, 74.59242, 73.8849, 73.15436, 73.78822, 74.9845,
  67.95179, 67.00564, 65.72301, 64.93632, 66.17059, 66.82233, 64.64048, 
    63.80264, 62.2719, 61.30988, 58.90459, 59.07368, 64.00903, 70.61009, 
    73.88804, 74.49326, 75.40926, 76.6992, 76.85645, 76.04742 ;
}
