netcdf tas_Amon_exAA01_historical_r1i1p1_198412-200511_box {
dimensions:
	lon = 20 ;
	bnds = 2 ;
	lat = 20 ;
	time = UNLIMITED ; // (4 currently)
variables:
	double lon(lon) ;
		lon:standard_name = "longitude" ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:axis = "X" ;
		lon:bounds = "lon_bnds" ;
	double lon_bnds(lon, bnds) ;
	double lat(lat) ;
		lat:standard_name = "latitude" ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:axis = "Y" ;
		lat:bounds = "lat_bnds" ;
	double lat_bnds(lat, bnds) ;
	double height ;
		height:standard_name = "height" ;
		height:long_name = "height" ;
		height:units = "m" ;
		height:positive = "up" ;
		height:axis = "Z" ;
	double time(time) ;
		time:standard_name = "time" ;
		time:long_name = "time" ;
		time:bounds = "time_bnds" ;
		time:units = "days since 1859-12-1 00:00:00" ;
		time:calendar = "360_day" ;
		time:axis = "T" ;
	double time_bnds(time, bnds) ;
	float tas(time, lat, lon) ;
		tas:standard_name = "air_temperature" ;
		tas:long_name = "Near-Surface Air Temperature" ;
		tas:units = "K" ;
		tas:coordinates = "height" ;
		tas:_FillValue = 1.e+20f ;
		tas:missing_value = 1.e+20f ;
		tas:comment = "near-surface (usually, 2 meter) air temperature." ;
		tas:original_name = "mo: m01s03i236" ;
		tas:cell_methods = "time: mean" ;
		tas:history = "2010-12-03T16:28:10Z altered by CMOR: Treated scalar dimension: \'height\'. 2010-12-03T16:28:10Z altered by CMOR: replaced missing value flag (-1.07374e+09) with standard missing value (1e+20)." ;
		tas:associated_files = "baseURL: http://cmip-pcmdi.llnl.gov/CMIP5/dataLocation gridspecFile: gridspec_atmos_fx_HadGEM2-ES_historical_r0i0p0.nc areacella: areacella_fx_HadGEM2-ES_historical_r0i0p0.nc" ;

// global attributes:
		:CDI = "Climate Data Interface version ?? (http://mpimet.mpg.de/cdi)" ;
		:Conventions = "CF-1.4" ;
		:history = "reset by cdo to create anonymous sample file" ;
		:source = "201707_compliance_checker_evaluation/work/p1.py" ;
		:institution = "CEDA" ;
		:institute_id = "CEDA" ;
		:experiment_id = "historical" ;
		:model_id = "exAA01" ;
		:forcing = "GHG, SA, Oz, LU, Sl, Vl, BC, OC, (GHG = CO2, N2O, CH4, CFCs)" ;
		:parent_experiment_id = "piControl" ;
		:parent_experiment_rip = "r1i1p1" ;
		:branch_time = 0. ;
		:contact = "none" ;
		:references = "Bellouin N. et al, (2007) Improved representation of aerosols for HadGEM2. Meteorological Office Hadley Centre, Technical Note 73, March 2007; Collins W.J.  et al, (2008) Evaluation of the HadGEM2 model. Meteorological Office Hadley Centre, Technical Note 74,; Johns T.C. et al, (2006) The new Hadley Centre climate model HadGEM1: Evaluation of coupled simulations. Journal of Climate, American Meteorological Society, Vol. 19, No. 7, pages 1327-1353.; Martin G.M. et al, (2006) The physical properties of the atmosphere in the new Hadley Centre Global Environmental Model, HadGEM1 - Part 1: Model description and global climatology. Journal of Climate, American Meteorological Society, Vol. 19, No.7, pages 1274-1301.; Ringer M.A. et al, (2006) The physical properties of the atmosphere in the new Hadley Centre Global Environmental Model, HadGEM1 - Part 2: Aspects of variability and regional climate. Journal of Climate, American Meteorological Society, Vol. 19, No. 7, pages 1302-1326." ;
		:initialization_method = 1 ;
		:physics_version = 1 ;
		:tracking_id = "c9bcc54c-aacb-4f5b-8ca0-23eaea5f6cbf" ;
		:mo_runid = "ajhoh" ;
		:product = "output" ;
		:experiment = "historical" ;
		:frequency = "mon" ;
		:creation_date = "2010-12-04T03:45:05Z" ;
		:project_id = "CMIP5" ;
		:table_id = "Table Amon (12 November 2010) 6e535ddfacb41fb7a252f4862fdc5766" ;
		:title = "Dummy file with known metadata errors" ;
		:parent_experiment = "pre-industrial control" ;
		:modeling_realm = "atmos" ;
		:realization = 1 ;
		:cmor_version = "2.5.0" ;
		:comment = "this is a sample file with known metadata errors" ;
		:CDO = "Climate Data Operators version 1.7.0 (http://mpimet.mpg.de/cdo)" ;
data:

 lon = 0, 1.875, 3.75, 5.625, 7.5, 9.375, 11.25, 13.125, 15, 16.875, 18.75, 
    20.625, 22.5, 24.375, 26.25, 28.125, 30, 31.875, 33.75, 35.625 ;

 lon_bnds =
  -0.9375, 0.9375,
  0.9375, 2.8125,
  2.8125, 4.6875,
  4.6875, 6.5625,
  6.5625, 8.4375,
  8.4375, 10.3125,
  10.3125, 12.1875,
  12.1875, 14.0625,
  14.0625, 15.9375,
  15.9375, 17.8125,
  17.8125, 19.6875,
  19.6875, 21.5625,
  21.5625, 23.4375,
  23.4375, 25.3125,
  25.3125, 27.1875,
  27.1875, 29.0625,
  29.0625, 30.9375,
  30.9375, 32.8125,
  32.8125, 34.6875,
  34.6875, 36.5625 ;

 lat = -90, -88.75, -87.5, -86.25, -85, -83.75, -82.5, -81.25, -80, -78.75, 
    -77.5, -76.25, -75, -73.75, -72.5, -71.25, -70, -68.75, -67.5, -66.25 ;

 lat_bnds =
  -90, -89.375,
  -89.375, -88.125,
  -88.125, -86.875,
  -86.875, -85.625,
  -85.625, -84.375,
  -84.375, -83.125,
  -83.125, -81.875,
  -81.875, -80.625,
  -80.625, -79.375,
  -79.375, -78.125,
  -78.125, -76.875,
  -76.875, -75.625,
  -75.625, -74.375,
  -74.375, -73.125,
  -73.125, -71.875,
  -71.875, -70.625,
  -70.625, -69.375,
  -69.375, -68.125,
  -68.125, -66.875,
  -66.875, -65.625 ;

 height = 1.5 ;

 time = 45015, 45045, 45075, 45105 ;

 time_bnds =
  45000, 45030,
  45030, 45060,
  45060, 45090,
  45090, 45120 ;

 tas =
  253.8957, 253.8957, 253.8957, 253.8957, 253.8957, 253.8957, 253.8957, 
    253.8957, 253.8957, 253.8957, 253.8957, 253.8957, 253.8957, 253.8957, 
    253.8957, 253.8957, 253.8957, 253.8957, 253.8957, 253.8957,
  254.8863, 254.8512, 254.8142, 254.7734, 254.733, 254.6923, 254.6522, 
    254.6129, 254.5679, 254.5226, 254.4824, 254.4396, 254.3892, 254.3432, 
    254.2979, 254.2485, 254.2046, 254.1514, 254.1034, 254.0593,
  255.8096, 255.717, 255.6244, 255.5383, 255.4445, 255.3527, 255.2679, 
    255.1891, 255.0984, 254.9954, 254.9048, 254.8129, 254.7127, 254.618, 
    254.5319, 254.4409, 254.3485, 254.2581, 254.1631, 254.0771,
  256.0389, 255.9312, 255.8245, 255.728, 255.6309, 255.5457, 255.4413, 
    255.3184, 255.2042, 255.0734, 254.9534, 254.8163, 254.6703, 254.5297, 
    254.3927, 254.2375, 254.08, 253.9139, 253.7524, 253.5972,
  256.4588, 256.3648, 256.2612, 256.1738, 256.0812, 255.9783, 255.8723, 
    255.7614, 255.668, 255.5665, 255.443, 255.2812, 255.1038, 254.8997, 
    254.6937, 254.4946, 254.2581, 254.0246, 253.7774, 253.5225,
  257.0399, 256.8353, 256.6606, 256.5067, 256.3653, 256.2534, 256.1422, 
    256.0252, 255.916, 255.8129, 255.673, 255.5003, 255.2998, 255.1024, 
    254.876, 254.6045, 254.3173, 253.9696, 253.5882, 253.1561,
  257.9153, 257.6675, 257.3967, 257.1689, 256.9535, 256.7954, 256.666, 
    256.5013, 256.3468, 256.123, 255.915, 255.7167, 255.4377, 255.1323, 
    254.8148, 254.4316, 254.0256, 253.5804, 252.9929, 252.4363,
  257.9331, 257.665, 257.3445, 257.0625, 256.7062, 256.4431, 256.2061, 
    256.0061, 255.6207, 255.332, 255.062, 254.7523, 254.3769, 254.0447, 
    253.6944, 253.2412, 252.7835, 252.384, 251.9109, 251.4422,
  257.1874, 256.9587, 256.6888, 256.3746, 256.046, 255.7283, 255.4235, 
    254.9815, 254.5919, 254.2514, 253.9832, 253.6145, 253.2034, 252.749, 
    252.3626, 252.009, 251.7645, 251.5203, 251.3032, 250.9642,
  256.2037, 255.9393, 255.5783, 255.1957, 254.7824, 254.4897, 254.1934, 
    253.6628, 253.259, 252.9206, 252.7485, 252.502, 252.088, 251.6741, 
    251.3402, 250.8157, 250.4076, 250.0022, 249.7506, 249.5449,
  255.1268, 254.5786, 254.1516, 253.7698, 253.1858, 252.6966, 252.3199, 
    251.8386, 251.5099, 251.1681, 251.0601, 250.7236, 250.3643, 250.0631, 
    249.9422, 249.6452, 249.2417, 248.8976, 248.7161, 248.7776,
  254.1077, 253.5508, 253.0239, 252.4781, 252.1757, 251.8209, 251.35, 
    250.9592, 250.6517, 250.566, 250.27, 249.8627, 249.6715, 249.6284, 
    249.3422, 249.1455, 248.8114, 248.5804, 248.3375, 248.0879,
  253.7905, 253.1672, 252.5542, 251.5536, 250.7817, 250.7576, 250.1553, 
    249.7548, 249.588, 249.4561, 249.4069, 249.0814, 248.8691, 248.879, 
    249.2659, 249.46, 249.7312, 249.832, 249.8823, 249.8456,
  255.3019, 254.5211, 253.4748, 252.3354, 251.2397, 250.8415, 250.2709, 
    250.2366, 250.6358, 250.7874, 251.1619, 251.4755, 251.6787, 252.0905, 
    252.6153, 252.8259, 253.0657, 252.998, 252.778, 252.4323,
  260.5541, 259.5001, 258.462, 257.2402, 256.2148, 255.6098, 255.5518, 
    256.0695, 256.6673, 257.3745, 258.2448, 258.7711, 259.1465, 259.4582, 
    259.4293, 259.3199, 258.965, 258.3267, 257.5023, 256.8258,
  263.2392, 266.6226, 264.1791, 263.6542, 263.0692, 262.7345, 262.5793, 
    262.7348, 263.0755, 263.492, 264.1844, 264.7742, 265.2902, 265.5424, 
    265.485, 265.1552, 264.704, 263.7125, 262.5222, 261.4669,
  267.7099, 264.8542, 262.525, 261.918, 261.1772, 260.7005, 260.4611, 
    260.5244, 260.6039, 260.9719, 261.6985, 262.8343, 264.0477, 265.207, 
    267.3621, 268.8454, 267.6806, 267.2822, 266.8436, 265.5074,
  270.9886, 270.799, 270.5464, 270.4376, 270.2759, 270.1794, 270.1461, 
    269.9896, 269.8635, 269.855, 269.8169, 269.7077, 269.6696, 269.7211, 
    269.8864, 270.0591, 270.1332, 270.4398, 268.3745, 270.0705,
  271.1502, 271.1333, 271.0531, 271.0195, 270.9529, 270.909, 270.9279, 
    270.8641, 270.7094, 270.6074, 270.5815, 270.5705, 270.5029, 270.4223, 
    270.4769, 270.5704, 270.6522, 270.6891, 270.5264, 270.4928,
  271.4689, 271.4795, 271.4694, 271.4124, 271.5194, 271.6699, 271.611, 
    271.4166, 271.3055, 271.2284, 271.3622, 271.5215, 271.3694, 271.1314, 
    271.0672, 271.0544, 271.0434, 270.9811, 271.0377, 271.0751,
  255.1298, 255.1298, 255.1298, 255.1298, 255.1298, 255.1298, 255.1298, 
    255.1298, 255.1298, 255.1298, 255.1298, 255.1298, 255.1298, 255.1298, 
    255.1298, 255.1298, 255.1298, 255.1298, 255.1298, 255.1298,
  256.0702, 256.0441, 256.0173, 255.9794, 255.9383, 255.8962, 255.8563, 
    255.8143, 255.7742, 255.7337, 255.6964, 255.6525, 255.6168, 255.5794, 
    255.5384, 255.4971, 255.4585, 255.4178, 255.3774, 255.3414,
  256.5861, 256.4936, 256.4001, 256.3, 256.202, 256.1039, 256.0073, 255.9111, 
    255.8162, 255.7245, 255.6329, 255.5449, 255.4592, 255.3768, 255.29, 
    255.2047, 255.116, 255.0331, 254.9561, 254.8792,
  256.8085, 256.7024, 256.5922, 256.4929, 256.3679, 256.2372, 256.0982, 
    255.9575, 255.8227, 255.6901, 255.5693, 255.4394, 255.3024, 255.1717, 
    255.0425, 254.9188, 254.801, 254.6907, 254.5761, 254.451,
  257.1705, 257.0664, 256.9461, 256.8162, 256.677, 256.5107, 256.3459, 
    256.1883, 256.0347, 255.8594, 255.7049, 255.5683, 255.4078, 255.2563, 
    255.0912, 254.947, 254.7784, 254.5565, 254.3195, 254.0529,
  257.9125, 257.7653, 257.6224, 257.4939, 257.3464, 257.1696, 257.0282, 
    256.8958, 256.6868, 256.5005, 256.3176, 256.1493, 255.9115, 255.6233, 
    255.3199, 255.0822, 254.7803, 254.4414, 254.0721, 253.6721,
  258.603, 258.4036, 258.2123, 258.0018, 257.8088, 257.6638, 257.5397, 
    257.3495, 257.0138, 256.8079, 256.5156, 256.1905, 255.8394, 255.4598, 
    255.073, 254.6547, 254.2486, 253.8193, 253.3667, 252.9525,
  258.6874, 258.3631, 258.0104, 257.7306, 257.4462, 257.1991, 256.9045, 
    256.5952, 256.3156, 256.0568, 255.7538, 255.4423, 255.028, 254.5895, 
    254.1352, 253.623, 253.19, 252.7488, 252.3159, 251.785,
  257.9451, 257.4951, 257.0094, 256.6019, 256.1658, 255.8101, 255.4535, 
    255.1583, 254.9027, 254.597, 254.2691, 254.0136, 253.7661, 253.326, 
    252.8902, 252.4348, 252.0179, 251.6652, 251.1953, 250.7842,
  256.726, 256.1789, 255.6609, 255.2247, 254.9212, 254.5435, 254.243, 
    253.9004, 253.6299, 253.2886, 252.9335, 252.6017, 252.2666, 251.9689, 
    251.631, 251.2446, 250.8299, 250.4365, 250.0527, 249.7795,
  255.6719, 255.1141, 254.7058, 254.3526, 254.0422, 253.7569, 253.4482, 
    252.9868, 252.6318, 252.3422, 252.0034, 251.6201, 251.207, 250.9886, 
    250.6462, 250.2842, 249.8857, 249.518, 249.1827, 249.0275,
  254.5312, 254.3859, 254.0833, 253.8868, 253.6992, 253.254, 252.9793, 
    252.3221, 251.8056, 251.4487, 251.113, 250.7289, 250.3364, 250.1087, 
    249.9086, 249.8035, 249.6194, 249.5302, 249.3466, 249.2321,
  254.2678, 254.4543, 253.8354, 253.2738, 252.5992, 251.9655, 251.4132, 
    251.0607, 250.7585, 250.4153, 250.2163, 250.1905, 250.085, 249.8831, 
    250.0695, 250.1832, 250.4637, 250.861, 251.1307, 250.9525,
  256.1225, 255.3829, 254.4167, 253.5271, 252.7159, 252.1154, 251.9995, 
    252.0336, 252.0616, 252.2949, 252.3173, 252.5419, 252.7813, 252.9797, 
    253.2718, 253.5884, 253.7912, 253.8839, 253.9329, 253.7155,
  262.2281, 261.2778, 260.1435, 258.9479, 258.0103, 257.4655, 257.2416, 
    257.3956, 257.975, 258.8102, 259.5148, 260.1454, 260.567, 260.9214, 
    261.0924, 260.7715, 260.2646, 259.5509, 258.6592, 257.9752,
  267.9958, 268.8691, 266.6969, 266.0466, 265.4966, 265.1514, 265.1292, 
    265.3512, 265.7553, 266.2941, 266.9086, 267.4498, 267.7458, 267.7839, 
    267.5278, 267.1245, 266.351, 265.1771, 264.116, 263.0379,
  270.9066, 269.6773, 268.1636, 268.0126, 267.8141, 267.7237, 267.6439, 
    267.3405, 267.3983, 267.7889, 268.5391, 269.3431, 270.0942, 270.7953, 
    271.4426, 270.8494, 270.0048, 269.3531, 268.4847, 267.6666,
  271.8805, 271.6719, 271.5803, 271.5757, 271.5287, 271.5042, 271.3915, 
    271.4197, 271.6654, 271.8115, 272.062, 272.3195, 272.4125, 272.1088, 
    271.6534, 271.3082, 271.2501, 271.1964, 270.9256, 271.2386,
  273.4199, 273.3135, 273.2726, 273.3115, 273.3795, 273.5544, 273.509, 
    273.546, 273.6889, 273.7955, 274.0051, 274.2161, 274.2348, 274.0494, 
    273.5314, 272.7152, 271.7384, 271.5627, 271.5319, 271.5754,
  274, 274.058, 274.033, 274.0444, 274.0758, 274.1851, 274.3469, 274.5355, 
    274.5868, 274.8436, 275.0149, 275.1531, 275.2716, 275.361, 275.3423, 
    275.3695, 274.9719, 274.5231, 274.3729, 274.387,
  237.6437, 237.6437, 237.6437, 237.6437, 237.6437, 237.6437, 237.6437, 
    237.6437, 237.6437, 237.6437, 237.6437, 237.6437, 237.6437, 237.6437, 
    237.6437, 237.6437, 237.6437, 237.6437, 237.6437, 237.6437,
  238.743, 238.6824, 238.6196, 238.5554, 238.4921, 238.4278, 238.3658, 
    238.3054, 238.2444, 238.1876, 238.1341, 238.0825, 238.0323, 237.9727, 
    237.902, 237.8354, 237.7701, 237.702, 237.6378, 237.5759,
  239.785, 239.6407, 239.508, 239.3806, 239.2574, 239.1378, 239.0203, 
    238.9044, 238.788, 238.675, 238.5613, 238.4467, 238.3201, 238.1971, 
    238.0751, 237.9634, 237.8575, 237.7659, 237.6867, 237.6099,
  239.9927, 239.72, 239.4728, 239.2651, 239.0907, 238.9384, 238.7941, 
    238.6631, 238.5472, 238.4302, 238.3306, 238.2518, 238.1686, 238.1328, 
    238.0731, 238.009, 237.9564, 237.9129, 237.8686, 237.827,
  239.4941, 239.1198, 238.7944, 238.5243, 238.3107, 238.1475, 238.0356, 
    237.9842, 237.9645, 237.9796, 238.0281, 238.1028, 238.181, 238.2534, 
    238.3415, 238.4291, 238.5229, 238.588, 238.6237, 238.6315,
  239.277, 238.8638, 238.5245, 238.2581, 238.042, 237.9051, 237.834, 237.844, 
    237.9493, 238.1036, 238.313, 238.5672, 238.8204, 239.023, 239.1996, 
    239.3376, 239.4261, 239.4963, 239.5338, 239.5324,
  240.754, 240.2042, 239.7162, 239.2987, 238.9354, 238.6949, 238.6111, 
    238.6588, 238.8235, 239.0387, 239.2411, 239.5103, 239.822, 240.0208, 
    240.1157, 240.1269, 240.0817, 240.0025, 239.8955, 239.7828,
  242.993, 242.3741, 241.7664, 241.2661, 240.8071, 240.4489, 240.2603, 
    240.2073, 240.2164, 240.2561, 240.3207, 240.4311, 240.5589, 240.6574, 
    240.6081, 240.423, 240.1769, 239.9135, 239.5992, 239.3024,
  243.7919, 243.1478, 242.6418, 242.1537, 241.6254, 241.2318, 241.0071, 
    240.8834, 240.7664, 240.6113, 240.4197, 240.1973, 239.9999, 239.8481, 
    239.7368, 239.5701, 239.3671, 239.2217, 238.9017, 238.4911,
  243.2235, 242.6554, 242.1376, 241.6008, 241.0803, 240.6381, 240.2623, 
    239.9129, 239.5857, 239.2352, 238.9017, 238.5565, 238.2745, 238.14, 
    238.1283, 238.1189, 238.1391, 238.3008, 238.1807, 237.8638,
  242.9629, 242.1118, 241.3088, 240.5363, 239.8444, 239.2254, 238.7054, 
    238.2982, 238.0679, 238.046, 237.9354, 237.8745, 237.6448, 237.6315, 
    237.8758, 238.1177, 238.1597, 238.0649, 237.8153, 237.5121,
  243.8341, 242.6528, 241.5894, 240.8221, 240.2201, 239.6199, 239.1804, 
    238.849, 238.7122, 238.9128, 238.8115, 238.77, 238.5808, 238.4879, 
    238.5271, 238.5385, 238.5458, 238.3839, 238.0513, 237.7957,
  244.5037, 243.5716, 242.8214, 242.1136, 241.466, 241.0117, 240.7707, 
    240.69, 240.576, 240.4342, 240.2, 240.0303, 239.9375, 240.1962, 240.5098, 
    240.6979, 240.7899, 240.8096, 240.6936, 240.4642,
  249.3917, 248.2343, 246.8369, 245.4589, 244.0834, 243.309, 242.9074, 
    242.9807, 243.1879, 243.3847, 243.759, 244.1953, 244.8182, 245.7213, 
    246.3414, 246.5147, 246.2399, 245.9369, 245.7458, 245.262,
  255.3487, 254.944, 254.3573, 253.3763, 252.3145, 251.7896, 251.5325, 
    251.606, 251.8073, 252.4291, 253.3038, 254.1705, 254.864, 255.3671, 
    255.376, 254.842, 253.8238, 253.1579, 252.4206, 251.7499,
  268.7853, 265.9279, 259.2272, 259.2481, 257.9906, 257.1597, 256.4932, 
    256.0712, 256.1399, 256.3804, 257.1355, 258.1739, 258.7934, 259.22, 
    259.189, 259.3498, 259.722, 258.9017, 258.2726, 257.5363,
  270.731, 270.6745, 270.0823, 270.1902, 270.1831, 270.1105, 269.8814, 
    269.7448, 269.8274, 269.6514, 269.2063, 269.6195, 270.5574, 271.0832, 
    271.6104, 269.2288, 262.8634, 263.0881, 262.5387, 263.0408,
  272.8409, 272.8153, 272.7986, 272.8828, 272.8585, 272.7995, 272.6748, 
    272.4968, 272.3519, 272.2767, 272.4254, 272.5291, 272.7039, 272.842, 
    272.9999, 272.8065, 272.0174, 271.9339, 269.0396, 270.2523,
  273.9214, 273.8524, 273.8751, 273.8733, 273.8888, 273.9305, 273.9496, 
    273.9783, 274.0259, 274.0758, 274.1891, 274.222, 274.3107, 274.2493, 
    274.2115, 274.1853, 273.9551, 273.5624, 272.4139, 272.7239,
  274.5945, 274.5676, 274.5829, 274.6223, 274.6725, 274.6693, 274.7372, 
    274.8182, 274.8999, 275.0428, 275.1896, 275.2988, 275.4001, 275.4349, 
    275.4156, 275.3698, 275.2905, 275.221, 275.08, 275.3055,
  225.4667, 225.4667, 225.4667, 225.4667, 225.4667, 225.4667, 225.4667, 
    225.4667, 225.4667, 225.4667, 225.4667, 225.4667, 225.4667, 225.4667, 
    225.4667, 225.4667, 225.4667, 225.4667, 225.4667, 225.4667,
  227.8345, 227.7933, 227.7769, 227.743, 227.6643, 227.6387, 227.5778, 
    227.4955, 227.4774, 227.4214, 227.3651, 227.3056, 227.26, 227.2109, 
    227.1406, 227.0619, 226.9874, 226.8987, 226.8193, 226.7214,
  228.4475, 228.2767, 228.1157, 227.9701, 227.8155, 227.6739, 227.532, 
    227.3646, 227.2098, 227.0737, 226.9465, 226.8413, 226.7396, 226.6331, 
    226.5215, 226.4059, 226.3004, 226.1901, 226.1117, 225.9977,
  228.2396, 227.9046, 227.5942, 227.3556, 227.1137, 226.8871, 226.6724, 
    226.441, 226.2399, 226.0197, 225.889, 225.7788, 225.6663, 225.5518, 
    225.4341, 225.2982, 225.1675, 225.0195, 224.8752, 224.7354,
  227.8485, 227.2631, 226.7054, 226.2238, 225.7838, 225.3958, 225.0609, 
    224.7991, 224.5892, 224.4418, 224.3613, 224.3162, 224.2972, 224.3083, 
    224.3276, 224.3554, 224.4175, 224.4614, 224.4688, 224.4172,
  227.9968, 227.3715, 226.8003, 226.2861, 225.8201, 225.4247, 225.0934, 
    224.8627, 224.7601, 224.7049, 224.7755, 224.8695, 224.9946, 225.1232, 
    225.2343, 225.3541, 225.4254, 225.4324, 225.3414, 225.16,
  230.8193, 230.0565, 229.3002, 228.639, 228.0554, 227.5392, 227.1521, 
    226.9153, 226.78, 226.7374, 226.7721, 226.9412, 227.1069, 227.0806, 
    227.0126, 226.853, 226.5705, 226.2214, 225.8149, 225.4116,
  234.6504, 233.6328, 232.6439, 231.7966, 231.0098, 230.4558, 230.1076, 
    229.8503, 229.7209, 229.6122, 229.5816, 229.6269, 229.5795, 229.3212, 
    228.8987, 228.3928, 227.773, 227.0875, 226.3359, 225.5882,
  235.9677, 234.6205, 233.542, 232.8254, 232.0941, 231.6868, 231.4791, 
    231.3983, 231.2437, 230.949, 230.5867, 230.0967, 229.5109, 228.9306, 
    228.5134, 228.2231, 227.9386, 227.5257, 226.7943, 225.7018,
  235.0765, 233.8231, 232.8812, 232.2006, 231.4675, 231.0563, 230.5436, 
    230.0438, 229.6308, 229.0967, 228.2716, 227.2642, 226.3489, 225.8165, 
    225.7942, 226.0416, 226.4263, 226.5784, 226.3923, 225.9131,
  234.8253, 233.5834, 232.2599, 231.0978, 229.9171, 228.7477, 227.8098, 
    227.1279, 226.9368, 227.2499, 227.0718, 226.7802, 226.256, 225.8359, 
    225.8615, 226.3299, 226.871, 227.1173, 226.9202, 226.3699,
  236.6445, 235.0801, 233.5166, 232.5095, 231.548, 230.6918, 229.8436, 
    229.1522, 228.9142, 229.5605, 229.4721, 229.154, 228.639, 228.3239, 
    228.1882, 228.201, 228.268, 227.866, 226.7495, 225.616,
  239.2803, 237.6818, 236.487, 235.8304, 235.2235, 234.7222, 233.9313, 
    233.1929, 232.7943, 232.8229, 232.4976, 232.3708, 232.4171, 232.3479, 
    232.2025, 232.2007, 232.0617, 231.7675, 231.3058, 230.5204,
  246.2079, 244.4246, 242.8799, 241.4382, 239.5933, 238.2484, 237.1281, 
    237.1926, 237.5523, 237.8558, 238.5897, 239.5037, 240.1818, 240.9458, 
    241.1359, 241.033, 240.6113, 240.3984, 240.3467, 239.7742,
  253.2656, 253.4681, 252.9084, 251.6967, 250.9933, 250.5025, 250.159, 
    249.95, 250.2073, 250.8469, 251.4736, 252.0855, 252.8499, 253.2347, 
    252.9275, 252.2346, 251.4437, 250.7217, 249.8398, 248.8594,
  266.3942, 263.319, 256.8201, 256.8017, 256.0684, 255.5054, 254.8774, 
    254.7573, 255.0338, 255.4644, 256.4164, 257.6874, 258.887, 259.1957, 
    259.592, 259.6138, 259.8025, 258.5019, 257.2841, 255.9526,
  271.3306, 271.2378, 270.5994, 270.6438, 270.2321, 270.0096, 269.6108, 
    269.1923, 268.6466, 268.2646, 268.4015, 269.0816, 269.9631, 270.5521, 
    270.6552, 268.7552, 264.7343, 264.4131, 263.2894, 263.7263,
  272.6682, 272.597, 272.528, 272.5237, 272.4387, 272.2984, 272.1606, 
    272.0995, 272.1699, 272.3126, 272.549, 272.9578, 273.3005, 273.3832, 
    273.3631, 273.129, 272.728, 272.3661, 270.2099, 271.3497,
  273.4522, 273.4752, 273.4828, 273.5323, 273.6131, 273.6738, 273.7267, 
    273.894, 274.105, 274.3543, 274.5021, 274.691, 274.7222, 274.7255, 
    274.705, 274.5984, 274.384, 274.0949, 272.5417, 272.8109,
  274.0247, 274.0922, 274.1573, 274.2942, 274.4514, 274.5958, 274.7155, 
    274.8887, 275.0151, 275.2092, 275.4171, 275.5736, 275.5822, 275.5487, 
    275.5028, 275.4037, 275.3592, 275.3887, 275.3625, 275.4565 ;
}
