netcdf hurs_Amon_bcc-csm1-1_decadal1981_r1i1p1_198201-199112_box {
dimensions:
	lon = 20 ;
	bnds = 2 ;
	lat = 20 ;
	time = UNLIMITED ; // (120 currently)
variables:
	double lon(lon) ;
		lon:standard_name = "longitude" ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:axis = "X" ;
		lon:bounds = "lon_bnds" ;
	double lon_bnds(lon, bnds) ;
	double lat(lat) ;
		lat:standard_name = "latitude" ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:axis = "Y" ;
		lat:bounds = "lat_bnds" ;
	double lat_bnds(lat, bnds) ;
	double height ;
		height:standard_name = "height" ;
		height:long_name = "height" ;
		height:units = "m" ;
		height:positive = "up" ;
		height:axis = "Z" ;
	double time(time) ;
		time:standard_name = "time" ;
		time:long_name = "time" ;
		time:bounds = "time_bnds" ;
		time:units = "days since 1982-1-1 00:00:00" ;
		time:calendar = "365_day" ;
		time:axis = "T" ;
	double time_bnds(time, bnds) ;
	float hurs(time, lat, lon) ;
		hurs:standard_name = "relative_humidity" ;
		hurs:long_name = "Near-Surface Relative Humidity" ;
		hurs:units = "%" ;
		hurs:grid_type = "gaussian" ;
		hurs:coordinates = "height" ;
		hurs:_FillValue = 1.e+20f ;
		hurs:missing_value = 1.e+20f ;
		hurs:comment = "This is the relative humidity with respect to liquid water for T> 0 C, and with respect to ice for T<0 C." ;
		hurs:original_name = "HURS" ;
		hurs:cell_methods = "time: mean (interval: 20 mintues)" ;
		hurs:history = "2012-08-15T07:31:53Z altered by CMOR: Treated scalar dimension: \'height\'." ;
		hurs:associated_files = "baseURL: http://cmip-pcmdi.llnl.gov/CMIP5/dataLocation gridspecFile: gridspec_atmos_fx_bcc-csm1-1_decadal1981_r0i0p0.nc areacella: areacella_fx_bcc-csm1-1_decadal1981_r0i0p0.nc" ;

// global attributes:
		:CDI = "Climate Data Interface version ?? (http://mpimet.mpg.de/cdi)" ;
		:Conventions = "CF-1.4" ;
		:history = "Tue Jul 18 21:56:00 2017: cdo selindexbox,1,20,1,20 hurs_Amon_bcc-csm1-1_decadal1981_r1i1p1_198201-199112.nc hurs_Amon_bcc-csm1-1_decadal1981_r1i1p1_198201-199112_box.nc\n",
			"Output from monthly mean data 2012-08-15T07:31:53Z CMOR rewrote data to comply with CF standards and CMIP5 requirements." ;
		:source = "bcc-csm1-1:atmosphere:  BCC_AGCM2.1 (T42L26); land: BCC_AVIM1.0;ocean: MOM4_L40 (tripolar, 1 lon x (1-1/3) lat, L40);sea ice: SIS (tripolar,1 lon x (1-1/3) lat)" ;
		:institution = "Beijing Climate Center(BCC),China Meteorological Administration,China" ;
		:institute_id = "BCC" ;
		:experiment_id = "decadal1981" ;
		:model_id = "dummy" ;
		:forcing = "Nat Ant GHG SD Oz Sl Vl SS Ds BC OC" ;
		:parent_experiment_id = "historical" ;
		:parent_experiment_rip = "r1i1p1" ;
		:branch_time = 1981. ;
		:contact = "Dr. Tongwen Wu (twwu@cma.gov.cn)" ;
		:comment = "The experiment starts from historical run at 1st Sep. 1981. With ocean initial conditions using the nudging method to observed temperature for the 1st Sep. 1981. The atmospheric and land compositions are prescribed as in the historical run (expt. 3.2) and the RCP4.5 scenario (expt. 4.1) beyond year 2005." ;
		:initialization_method = 1 ;
		:physics_version = 1 ;
		:tracking_id = "37994f26-9f35-4e36-b539-8c9cdfa36487" ;
		:product = "output" ;
		:experiment = "10- or 30-year run initialized in year 1981" ;
		:frequency = "mon" ;
		:creation_date = "2012-08-15T07:31:54Z" ;
		:project_id = "CMIP5" ;
		:table_id = "Table Amon (11 April 2011) 1cfdc7322cf2f4a32614826fab42c1ab" ;
		:title = "bcc-csm1-1 model output prepared for CMIP5 10- or 30-year run initialized in year 1981" ;
		:parent_experiment = "historical" ;
		:modeling_realm = "atmos" ;
		:realization = 1 ;
		:cmor_version = "2.5.6" ;
		:CDO = "Climate Data Operators version 1.7.0 (http://mpimet.mpg.de/cdo)" ;
data:

 lon = 0, 2.8125, 5.625, 8.4375, 11.25, 14.0625, 16.875, 19.6875, 22.5, 
    25.3125, 28.125, 30.9375, 33.75, 36.5625, 39.375, 42.1875, 45, 47.8125, 
    50.625, 53.4375 ;

 lon_bnds =
  -1.40625, 1.40625,
  1.40625, 4.21875,
  4.21875, 7.03125,
  7.03125, 9.84375,
  9.84375, 12.65625,
  12.65625, 15.46875,
  15.46875, 18.28125,
  18.28125, 21.09375,
  21.09375, 23.90625,
  23.90625, 26.71875,
  26.71875, 29.53125,
  29.53125, 32.34375,
  32.34375, 35.15625,
  35.15625, 37.96875,
  37.96875, 40.78125,
  40.78125, 43.59375,
  43.59375, 46.40625,
  46.40625, 49.21875,
  49.21875, 52.03125,
  52.03125, 54.84375 ;

 lat = -87.8637988392326, -85.0965269883174, -82.3129129478863, 
    -79.5256065726594, -76.7368996803683, -73.9475151539897, 
    -71.1577520115873, -68.3677561083132, -65.5776070108278, 
    -62.7873517989631, -59.9970201084913, -57.2066315276432, 
    -54.4161995260862, -51.6257336749383, -48.8352409662506, 
    -46.0447266311017, -43.2541946653509, -40.463648178115, 
    -37.6730896290453, -34.8825209937735 ;

 lat_bnds =
  -87.8637988392326, -86.480162913775,
  -86.480162913775, -83.7047199681018,
  -83.7047199681018, -80.9192597602729,
  -80.9192597602729, -78.1312531265139,
  -78.1312531265139, -75.342207417179,
  -75.342207417179, -72.5526335827885,
  -72.5526335827885, -69.7627540599503,
  -69.7627540599503, -66.9726815595705,
  -66.9726815595705, -64.1824794048954,
  -64.1824794048954, -61.3921859537272,
  -61.3921859537272, -58.6018258180673,
  -58.6018258180673, -55.8114155268647,
  -55.8114155268647, -53.0209666005122,
  -53.0209666005122, -50.2304873205944,
  -50.2304873205944, -47.4399837986761,
  -47.4399837986761, -44.6494606482263,
  -44.6494606482263, -41.858921421733,
  -41.858921421733, -39.0683689035802,
  -39.0683689035802, -36.2778053114094,
  -36.2778053114094, -33.4872324377587 ;

 height = 2 ;

 time = 15.5, 45, 74.5, 105, 135.5, 166, 196.5, 227.5, 258, 288.5, 319, 
    349.5, 380.5, 410, 439.5, 470, 500.5, 531, 561.5, 592.5, 623, 653.5, 684, 
    714.5, 745.5, 775, 804.5, 835, 865.5, 896, 926.5, 957.5, 988, 1018.5, 
    1049, 1079.5, 1110.5, 1140, 1169.5, 1200, 1230.5, 1261, 1291.5, 1322.5, 
    1353, 1383.5, 1414, 1444.5, 1475.5, 1505, 1534.5, 1565, 1595.5, 1626, 
    1656.5, 1687.5, 1718, 1748.5, 1779, 1809.5, 1840.5, 1870, 1899.5, 1930, 
    1960.5, 1991, 2021.5, 2052.5, 2083, 2113.5, 2144, 2174.5, 2205.5, 2235, 
    2264.5, 2295, 2325.5, 2356, 2386.5, 2417.5, 2448, 2478.5, 2509, 2539.5, 
    2570.5, 2600, 2629.5, 2660, 2690.5, 2721, 2751.5, 2782.5, 2813, 2843.5, 
    2874, 2904.5, 2935.5, 2965, 2994.5, 3025, 3055.5, 3086, 3116.5, 3147.5, 
    3178, 3208.5, 3239, 3269.5, 3300.5, 3330, 3359.5, 3390, 3420.5, 3451, 
    3481.5, 3512.5, 3543, 3573.5, 3604, 3634.5 ;

 time_bnds =
  0, 31,
  31, 59,
  59, 90,
  90, 120,
  120, 151,
  151, 181,
  181, 212,
  212, 243,
  243, 273,
  273, 304,
  304, 334,
  334, 365,
  365, 396,
  396, 424,
  424, 455,
  455, 485,
  485, 516,
  516, 546,
  546, 577,
  577, 608,
  608, 638,
  638, 669,
  669, 699,
  699, 730,
  730, 761,
  761, 789,
  789, 820,
  820, 850,
  850, 881,
  881, 911,
  911, 942,
  942, 973,
  973, 1003,
  1003, 1034,
  1034, 1064,
  1064, 1095,
  1095, 1126,
  1126, 1154,
  1154, 1185,
  1185, 1215,
  1215, 1246,
  1246, 1276,
  1276, 1307,
  1307, 1338,
  1338, 1368,
  1368, 1399,
  1399, 1429,
  1429, 1460,
  1460, 1491,
  1491, 1519,
  1519, 1550,
  1550, 1580,
  1580, 1611,
  1611, 1641,
  1641, 1672,
  1672, 1703,
  1703, 1733,
  1733, 1764,
  1764, 1794,
  1794, 1825,
  1825, 1856,
  1856, 1884,
  1884, 1915,
  1915, 1945,
  1945, 1976,
  1976, 2006,
  2006, 2037,
  2037, 2068,
  2068, 2098,
  2098, 2129,
  2129, 2159,
  2159, 2190,
  2190, 2221,
  2221, 2249,
  2249, 2280,
  2280, 2310,
  2310, 2341,
  2341, 2371,
  2371, 2402,
  2402, 2433,
  2433, 2463,
  2463, 2494,
  2494, 2524,
  2524, 2555,
  2555, 2586,
  2586, 2614,
  2614, 2645,
  2645, 2675,
  2675, 2706,
  2706, 2736,
  2736, 2767,
  2767, 2798,
  2798, 2828,
  2828, 2859,
  2859, 2889,
  2889, 2920,
  2920, 2951,
  2951, 2979,
  2979, 3010,
  3010, 3040,
  3040, 3071,
  3071, 3101,
  3101, 3132,
  3132, 3163,
  3163, 3193,
  3193, 3224,
  3224, 3254,
  3254, 3285,
  3285, 3316,
  3316, 3344,
  3344, 3375,
  3375, 3405,
  3405, 3436,
  3436, 3466,
  3466, 3497,
  3497, 3528,
  3528, 3558,
  3558, 3589,
  3589, 3619,
  3619, 3650 ;

 hurs =
  93.4809, 93.74128, 93.9556, 94.03909, 94.47622, 94.65362, 94.82246, 
    95.1601, 93.7446, 94.10422, 94.16572, 94.11856, 94.13337, 94.49639, 
    94.70043, 94.81069, 93.98279, 94.30159, 94.16895, 94.13051,
  88.7273, 89.54988, 90.32349, 91.12242, 92.00128, 92.69608, 93.63831, 
    94.38155, 91.08723, 91.9362, 92.52862, 93.34216, 93.92194, 94.5956, 
    94.90078, 95.31381, 93.43739, 94.07809, 94.69255, 95.03079,
  83.48702, 84.99387, 86.29594, 87.70504, 88.8302, 89.77134, 91.012, 
    92.43107, 88.70104, 89.85878, 90.94014, 92.18761, 92.81371, 93.41303, 
    93.52509, 94.11451, 92.28455, 92.71619, 93.31631, 93.52835,
  84.69096, 86.19128, 87.67854, 89.19056, 90.50443, 91.71695, 92.53498, 
    93.33336, 90.69014, 91.27824, 91.97832, 92.61449, 93.1025, 93.40945, 
    93.54196, 93.37686, 93.75618, 93.67755, 93.39366, 93.51973,
  83.67885, 86.10898, 88.38322, 90.29052, 91.65009, 92.62195, 93.09725, 
    93.88835, 91.5418, 91.3267, 91.20734, 91.85376, 92.48512, 92.65701, 
    92.91588, 92.77927, 96.84536, 96.78885, 96.07845, 95.499,
  82.51562, 84.88831, 86.97651, 88.77648, 89.76414, 90.14468, 90.25821, 
    90.01252, 85.492, 85.72311, 86.30702, 87.01633, 88.00871, 89.5621, 
    91.02483, 92.61087, 98.50533, 98.64861, 98.5509, 98.17497,
  89.68507, 86.78841, 86.6087, 86.84266, 86.71143, 86.51164, 86.33993, 
    85.93306, 77.86455, 77.40113, 77.35551, 79.10056, 81.01414, 85.01857, 
    84.12335, 87.63353, 94.95633, 96.56116, 97.33598, 97.23394,
  93.43623, 92.90776, 91.67722, 90.48186, 89.21488, 88.15541, 87.04222, 
    85.63926, 77.28253, 75.64349, 75.49283, 78.94083, 78.86671, 79.91819, 
    70.37437, 74.3143, 78.09537, 93.66832, 94.12508, 95.66349,
  87.42145, 88.93051, 90.46446, 91.42157, 91.6532, 91.33952, 90.35046, 
    88.95781, 84.75066, 83.16238, 82.43893, 82.44582, 83.63319, 84.69102, 
    85.57793, 86.90664, 88.29635, 88.45477, 91.93355, 94.33942,
  84.33488, 86.3585, 88.88643, 91.39141, 92.21031, 91.9331, 91.31547, 
    90.97707, 90.83997, 90.39748, 90.02382, 89.0844, 88.53478, 88.39187, 
    88.94681, 89.19878, 89.81826, 91.08138, 92.13571, 92.45863,
  81.94168, 82.978, 84.72486, 87.94966, 90.65647, 91.54073, 91.38587, 
    91.50724, 92.07696, 92.36807, 92.84383, 92.41033, 91.17633, 90.46159, 
    90.12606, 89.69244, 89.76153, 89.78741, 90.41199, 91.27546,
  82.42509, 82.66344, 83.24526, 85.00698, 86.61463, 86.95371, 86.59507, 
    87.69249, 90.12206, 91.88249, 92.80717, 92.99869, 92.13709, 91.56483, 
    91.09361, 89.98956, 89.55358, 89.58495, 89.884, 90.68936,
  85.83164, 85.98697, 86.30321, 86.7794, 86.6998, 84.66866, 81.7151, 
    81.01419, 83.48742, 86.76139, 89.18749, 90.869, 91.45655, 91.09351, 
    91.39294, 91.30672, 90.09115, 88.65224, 88.784, 89.37923,
  82.37218, 83.16448, 83.78975, 84.20922, 83.2514, 81.95366, 81.78837, 
    82.77064, 84.525, 86.61893, 87.79867, 88.67591, 89.51363, 90.13094, 
    91.13078, 91.47941, 89.81043, 88.1453, 87.87795, 89.09147,
  75.86752, 75.09309, 75.2433, 75.39053, 75.22278, 76.72486, 80.25311, 
    83.74046, 86.40416, 87.6395, 88.04431, 88.57058, 89.66587, 90.52764, 
    90.9056, 91.11395, 90.21503, 89.09438, 89.44652, 90.82539,
  73.35105, 72.47985, 72.89262, 74.36884, 76.2441, 78.83097, 82.01714, 
    84.33385, 86.53508, 88.42753, 89.38844, 89.757, 90.1792, 90.89043, 
    91.0164, 90.70487, 89.87632, 89.47755, 90.27154, 90.51128,
  76.63313, 77.2861, 78.97208, 80.56419, 81.63042, 82.18461, 82.20987, 
    82.44176, 84.14093, 86.33018, 88.35344, 89.31207, 89.28953, 89.42931, 
    89.32444, 88.2574, 86.47741, 85.4045, 84.93102, 84.50637,
  83.00284, 82.76088, 82.8689, 81.82735, 80.72785, 79.71549, 79.37939, 
    78.76436, 74.75816, 73.10941, 74.78475, 78.0412, 80.88372, 82.72076, 
    84.10639, 84.26265, 82.52142, 79.37403, 77.83792, 78.10139,
  81.83013, 80.74139, 79.26865, 77.1935, 75.92776, 76.23385, 75.38225, 
    69.07002, 63.52311, 61.11913, 61.72075, 65.10432, 69.99793, 74.59365, 
    78.36984, 79.33351, 78.0505, 77.30078, 78.44856, 80.42095,
  73.47881, 72.02462, 70.44322, 69.69109, 69.98117, 70.39768, 67.90502, 
    63.09711, 60.43573, 58.8373, 59.27411, 63.01844, 70.89108, 76.50346, 
    78.50382, 78.2642, 78.4737, 79.86833, 81.52776, 82.52912,
  91.05083, 91.30476, 91.53485, 92.02209, 92.18385, 92.56113, 92.62751, 
    93.08926, 91.88125, 92.40703, 92.5981, 92.64035, 92.99768, 92.64845, 
    93.51599, 93.89808, 92.04053, 93.13046, 92.65516, 93.22881,
  86.96413, 87.80626, 88.72099, 89.57648, 90.3923, 91.21534, 92.04106, 
    92.90271, 89.44534, 90.34664, 91.18976, 92.07103, 92.96951, 93.7209, 
    94.42259, 95.10692, 93.32484, 94.06727, 94.6227, 94.98904,
  85.80513, 87.10407, 88.54015, 89.99532, 91.11778, 92.29962, 93.42702, 
    94.41877, 90.26347, 91.3447, 92.29098, 93.48471, 94.67207, 95.65806, 
    96.47842, 97.24012, 95.63651, 96.28072, 96.89655, 97.20786,
  85.95926, 87.22572, 88.69738, 90.30405, 91.83503, 92.93233, 94.13572, 
    95.26557, 93.02795, 94.30644, 95.31511, 95.90936, 96.54295, 97.02541, 
    97.50476, 97.7431, 98.66412, 98.55714, 98.53976, 97.77951,
  84.73331, 86.33834, 88.74374, 90.77811, 92.45103, 93.38811, 94.29533, 
    95.24791, 94.00957, 94.55647, 94.90408, 95.08174, 95.35646, 96.20399, 
    96.47029, 96.29651, 99.09619, 98.84468, 98.37006, 97.46123,
  84.39301, 86.8561, 88.84941, 90.42979, 91.79298, 92.48118, 92.73416, 
    92.78191, 88.05251, 88.12733, 88.48933, 88.75777, 89.77502, 90.84673, 
    91.97835, 93.42875, 98.78717, 98.84388, 98.49764, 98.00574,
  88.28484, 85.12112, 84.33315, 84.39015, 84.37801, 84.40788, 84.34162, 
    84.17943, 76.47164, 75.87708, 75.25665, 74.02428, 76.02343, 84.70475, 
    85.37189, 84.09641, 92.42211, 95.36664, 96.6904, 97.2202,
  70.56541, 68.4983, 67.41721, 66.8833, 67.7931, 69.21661, 69.8529, 69.42115, 
    63.17681, 62.5233, 62.89027, 67.26984, 66.06211, 65.23525, 55.66279, 
    58.71144, 67.86268, 87.54339, 86.85458, 88.93345,
  68.84487, 68.51212, 69.35588, 71.91167, 74.11705, 75.94108, 76.46138, 
    75.37688, 71.65511, 70.68373, 70.22173, 70.43938, 71.64607, 72.97045, 
    74.19555, 75.15436, 74.11209, 71.4112, 75.65611, 78.24518,
  76.204, 75.76051, 76.30462, 78.38274, 80.0094, 80.87751, 81.61044, 
    81.53532, 81.66994, 81.50655, 81.2676, 81.04417, 81.54856, 82.12254, 
    81.42691, 81.53082, 82.43788, 82.96621, 83.54175, 83.96078,
  80.23288, 79.93113, 79.55199, 80.25504, 81.74779, 82.56519, 82.99827, 
    83.67518, 84.84621, 85.20068, 86.04611, 86.85261, 87.18818, 86.70637, 
    85.09091, 83.79376, 83.47128, 83.66501, 84.92827, 87.11862,
  80.3205, 80.81688, 80.38798, 80.2877, 80.36696, 80.49259, 80.68171, 
    81.90107, 84.04259, 86.0901, 87.90427, 89.13175, 89.38041, 88.99027, 
    87.82668, 86.39554, 85.45226, 85.01891, 85.1569, 85.85855,
  82.61204, 84.35664, 84.58595, 83.7952, 83.19865, 82.12931, 80.47408, 
    80.31496, 81.63389, 84.10897, 86.23838, 88.20938, 89.64275, 90.14081, 
    90.22598, 89.43638, 87.71576, 85.99191, 85.64497, 86.32988,
  77.52943, 80.00568, 81.99464, 82.82799, 82.7672, 81.90527, 81.63331, 
    82.93295, 84.85116, 86.85659, 88.73515, 90.06676, 91.00152, 91.6852, 
    92.33061, 92.27951, 91.1763, 90.12089, 90.0131, 90.05972,
  70.85555, 71.13307, 72.69428, 75.08057, 76.58379, 77.37475, 79.43566, 
    82.78063, 85.86054, 88.28426, 90.07277, 91.17024, 91.87083, 91.45269, 
    90.72025, 90.61872, 90.62669, 90.56753, 90.9033, 91.29102,
  67.00684, 67.09906, 68.57079, 71.75898, 74.98229, 77.92363, 81.4397, 
    83.80692, 85.61021, 87.91116, 89.82823, 90.51535, 90.31052, 89.72369, 
    89.45454, 89.80968, 89.86005, 89.7135, 90.07793, 89.7205,
  67.42973, 69.64367, 73.03672, 76.33788, 78.47476, 80.10015, 81.0109, 
    81.44915, 82.62988, 84.73471, 86.24037, 86.77477, 86.97071, 87.5002, 
    87.86768, 87.51228, 86.24092, 84.8092, 83.44328, 81.98793,
  71.84314, 73.90975, 76.41698, 77.60235, 77.50567, 77.15674, 76.7172, 
    76.34422, 73.36298, 72.05531, 73.5601, 76.21287, 79.43002, 81.82706, 
    82.31962, 81.0184, 78.15611, 74.86246, 73.23536, 72.86601,
  72.87029, 73.06731, 73.01364, 72.42223, 71.79234, 72.95309, 72.38346, 
    67.12737, 64.14597, 63.28709, 64.52564, 67.76785, 72.1254, 74.02386, 
    73.94988, 72.74982, 70.37342, 69.23614, 70.56975, 72.32249,
  66.57248, 65.85196, 64.97097, 64.76868, 66.37942, 68.13031, 66.52633, 
    63.15863, 64.16334, 65.31944, 65.01894, 65.8837, 69.25704, 71.14582, 
    70.45712, 69.66892, 70.43227, 72.44795, 74.49334, 76.20102,
  92.22964, 92.43774, 92.63062, 92.8927, 93.19102, 93.51788, 93.97072, 
    94.11161, 92.57564, 92.95654, 92.68084, 92.93453, 92.90622, 93.64265, 
    93.20396, 93.64107, 92.85706, 93.42496, 93.58959, 94.07526,
  86.53026, 87.48244, 88.50666, 89.69047, 90.90907, 91.94442, 92.98344, 
    94.28337, 91.34309, 92.40143, 93.23909, 93.97713, 94.6262, 95.10246, 
    95.59241, 96.23475, 94.76723, 95.52543, 96.14085, 96.77498,
  86.57798, 88.27718, 90.18165, 92.02053, 93.36674, 94.7112, 95.64027, 
    96.24773, 92.06914, 93.2021, 94.23994, 95.49935, 96.77421, 97.63377, 
    97.98104, 98.39999, 97.01608, 97.34422, 97.65852, 98.02956,
  85.57472, 87.42229, 89.42072, 91.31242, 92.87572, 94.0182, 94.81004, 
    95.25046, 92.9412, 93.63285, 94.24619, 94.66399, 95.5916, 96.98648, 
    97.69051, 97.93504, 98.9244, 99.30836, 99.28754, 99.01913,
  79.8897, 81.06566, 83.05697, 84.85406, 86.71394, 88.3033, 89.21417, 
    90.49871, 89.98582, 90.96175, 90.5547, 91.20617, 91.58131, 92.33372, 
    92.52147, 92.46666, 95.38915, 95.59892, 95.88333, 95.71642,
  81.32919, 83.57585, 85.60041, 87.10515, 87.96142, 88.2849, 88.83413, 
    89.01068, 84.51334, 84.6098, 85.05444, 85.95848, 86.76998, 87.46896, 
    87.9019, 88.61512, 94.58236, 95.06998, 95.14769, 94.7646,
  88.07307, 86.59868, 86.58923, 85.98232, 87.31383, 89.03308, 87.69571, 
    86.28378, 78.07515, 77.42992, 76.50029, 75.31867, 77.60992, 84.57999, 
    88.4496, 83.90228, 90.68993, 92.63293, 93.92556, 94.3019,
  66.82751, 64.60086, 62.82958, 61.60794, 63.41624, 65.40393, 63.58063, 
    61.02935, 54.88851, 52.43182, 52.38718, 59.72296, 63.81407, 71.09298, 
    73.98959, 77.97992, 85.19641, 87.71232, 85.54469, 85.85326,
  73.13551, 71.02815, 69.26849, 68.40961, 68.70718, 70.467, 72.87477, 
    74.51218, 72.79417, 72.56232, 72.75586, 73.20984, 73.98312, 74.24403, 
    72.93912, 70.91954, 68.17037, 66.61717, 71.47506, 76.72422,
  79.34602, 78.66451, 78.3548, 77.70069, 76.63519, 76.07726, 76.30894, 
    76.85977, 77.66917, 78.23744, 78.81143, 79.5592, 80.23734, 80.9165, 
    81.75278, 81.83458, 81.53395, 81.31597, 81.78459, 81.8632,
  82.1837, 81.05145, 80.16758, 79.96313, 79.35477, 78.85178, 79.16402, 
    79.59003, 80.19248, 80.37486, 80.93359, 81.53082, 82.25062, 83.12988, 
    83.54334, 83.05065, 82.54458, 82.45341, 83.38203, 85.05447,
  82.27977, 81.84331, 81.39489, 81.61255, 81.11818, 80.31812, 79.75488, 
    80.21078, 81.15015, 82.00865, 82.57651, 82.95551, 83.45312, 84.68269, 
    85.90909, 85.93105, 85.15443, 84.02096, 83.69626, 84.02985,
  83.19819, 84.77756, 85.29516, 85.23341, 84.3204, 81.84599, 78.9753, 
    78.56066, 80.26664, 82.85178, 84.57373, 85.59086, 86.2681, 87.16847, 
    88.62134, 89.42458, 88.9723, 87.42092, 86.10884, 85.40966,
  77.55661, 78.20733, 78.97232, 78.85659, 77.29427, 75.32452, 73.60342, 
    73.67761, 76.62664, 80.55087, 83.18075, 85.25797, 87.23463, 89.3175, 
    91.49753, 91.87869, 91.04417, 90.20111, 89.73278, 89.18158,
  72.69135, 71.18095, 70.91507, 71.17534, 70.98412, 71.0764, 71.73852, 
    74.35057, 78.77151, 82.15887, 84.43987, 86.56584, 88.47732, 90.17076, 
    91.45909, 91.71172, 91.01821, 90.18664, 90.21486, 90.02959,
  71.88069, 70.26759, 69.84135, 70.97539, 72.88988, 75.61446, 78.73995, 
    81.53966, 83.13571, 84.78057, 86.86706, 88.44273, 89.37089, 89.90425, 
    89.52814, 88.78856, 87.91721, 86.92907, 87.05277, 86.4493,
  75.1648, 75.33139, 76.83544, 78.9208, 80.75966, 81.75249, 81.45548, 
    80.67786, 81.05466, 83.27165, 85.56857, 86.81513, 87.19731, 87.20964, 
    85.99469, 84.66291, 83.5312, 82.70512, 82.69513, 82.53698,
  80.13885, 80.93002, 82.51959, 82.78947, 81.56464, 79.74812, 78.35667, 
    76.45396, 71.82506, 70.24403, 72.7714, 76.51721, 79.09177, 80.22096, 
    81.24654, 81.64393, 80.49542, 79.13195, 78.72643, 78.86671,
  78.32669, 78.63792, 78.58054, 76.83755, 75.471, 75.81986, 74.33036, 
    67.22467, 61.09481, 59.61237, 61.09739, 64.24065, 68.30055, 72.31342, 
    76.53555, 78.25968, 77.88239, 77.30264, 77.3987, 77.07419,
  68.94539, 68.68242, 67.90125, 67.52906, 68.38454, 68.82463, 66.44341, 
    64.24481, 64.48137, 66.51134, 66.76366, 67.10056, 71.16967, 76.8642, 
    79.77894, 78.94858, 78.6658, 79.55561, 79.34438, 78.17169,
  92.54141, 93.03654, 93.52762, 93.84403, 94.29354, 94.51123, 94.85713, 
    95.37252, 93.90202, 94.31615, 94.88012, 95.2742, 95.43367, 95.5916, 
    95.6601, 95.76815, 94.76352, 94.81911, 95.11162, 94.88686,
  88.01664, 89.33185, 90.5452, 91.72334, 93.03945, 94.02189, 94.6624, 
    95.15916, 91.48368, 92.13939, 92.6049, 93.2338, 94.24551, 95.44672, 
    96.71396, 97.30254, 96.08929, 97.30815, 98.098, 98.56557,
  90.94303, 92.52785, 93.59134, 94.15833, 94.02104, 94.04562, 94.29615, 
    95.22523, 92.14843, 93.13724, 94.34363, 95.3501, 95.84255, 96.49215, 
    97.14639, 97.7093, 96.85003, 96.86707, 98.12727, 98.75555,
  88.27318, 90.09724, 90.99214, 92.27362, 93.60272, 94.15263, 94.1814, 
    93.75691, 92.58743, 94.21455, 95.44579, 95.48254, 97.53008, 98.88947, 
    99.46278, 99.73093, 99.77509, 99.8382, 99.89862, 99.71155,
  87.89031, 90.40994, 91.82758, 92.53615, 90.4079, 89.04392, 86.26049, 
    84.59306, 84.01423, 84.81204, 87.06075, 90.74068, 92.94947, 94.75008, 
    96.19665, 97.18544, 98.77139, 98.6069, 98.57997, 98.00607,
  83.8903, 84.92136, 85.39373, 85.37511, 84.69858, 83.02608, 82.80133, 
    82.95575, 79.49889, 80.70763, 82.39478, 84.50827, 86.53953, 88.32211, 
    89.75426, 90.74025, 97.06171, 97.45334, 97.07273, 96.55278,
  90.88854, 89.76771, 89.11231, 88.62409, 87.96299, 88.64448, 89.22742, 
    89.59662, 83.00499, 84.28205, 85.38667, 75.99948, 78.06296, 86.1804, 
    91.22605, 85.66981, 91.63414, 93.50183, 94.56201, 95.41918,
  68.94415, 66.33955, 64.29183, 65.86238, 68.57698, 72.97327, 75.46369, 
    75.94781, 70.16953, 71.42984, 75.55386, 78.06153, 82.2213, 89.04475, 
    92.60138, 93.229, 94.92187, 93.98281, 90.93874, 89.7681,
  71.95364, 69.37602, 67.37003, 65.48115, 64.44978, 64.15454, 64.02914, 
    64.00714, 62.10726, 62.3767, 63.09856, 64.20993, 65.98297, 68.32056, 
    69.56511, 70.84837, 74.83064, 81.55328, 86.19711, 88.44236,
  80.79776, 81.13727, 80.99896, 80.06807, 78.51117, 76.4956, 74.8095, 
    73.18134, 72.48692, 72.22964, 72.51437, 73.08861, 73.94782, 75.33536, 
    76.24101, 76.79229, 77.74096, 77.86268, 77.6832, 76.9064,
  82.41901, 82.753, 82.95709, 83.02888, 82.5001, 81.62798, 80.52926, 
    79.42319, 79.03169, 78.65395, 78.60709, 78.77505, 79.4987, 80.38777, 
    80.64737, 80.33028, 80.24097, 79.32241, 78.44655, 78.81319,
  82.85352, 83.37037, 83.26756, 83.29868, 82.87095, 81.83881, 81.79357, 
    83.27275, 85.26991, 85.91756, 85.69547, 85.26593, 85.25497, 85.41699, 
    85.35724, 84.64681, 83.86331, 82.14967, 80.87762, 80.50623,
  83.38592, 85.35951, 86.53141, 86.30074, 85.66002, 84.33922, 81.94282, 
    80.93518, 81.83748, 83.32011, 84.69791, 86.03635, 87.139, 87.7773, 
    88.77158, 89.18918, 88.49197, 86.56252, 84.66927, 82.93718,
  75.79934, 76.75446, 77.52898, 77.5277, 76.99945, 76.20707, 75.2501, 
    74.26753, 74.8577, 77.57658, 80.82764, 84.20567, 87.21058, 89.12047, 
    90.78375, 91.23209, 90.35426, 89.3278, 88.5433, 86.92542,
  69.21698, 68.35692, 68.80516, 69.58924, 70.05959, 70.75885, 71.75528, 
    73.23194, 77.27584, 82.16837, 86.12025, 88.95671, 90.60925, 90.88049, 
    90.78745, 90.44984, 89.46867, 88.44221, 88.83672, 89.24079,
  68.50562, 68.10552, 68.59997, 70.33549, 72.60332, 75.29845, 78.04709, 
    80.88697, 83.91629, 86.45277, 88.43858, 89.40572, 89.91223, 90.19718, 
    90.01281, 89.71179, 89.20315, 88.67767, 89.69603, 89.97243,
  71.52088, 73.22936, 75.69386, 78.65891, 81.17647, 82.8969, 83.16904, 
    82.24049, 81.93842, 83.45264, 86.2891, 87.97657, 88.5819, 88.9337, 
    88.85368, 88.32925, 87.61467, 86.53557, 86.01635, 85.59343,
  75.79662, 78.00786, 80.5469, 81.59884, 80.70174, 78.97758, 77.41759, 
    74.14724, 69.33091, 69.06882, 72.36685, 76.35325, 79.35719, 81.87857, 
    83.53662, 83.43586, 81.40395, 78.64791, 77.64761, 78.19087,
  75.40871, 75.86194, 75.55762, 73.83998, 72.1325, 71.50379, 69.34479, 
    62.2871, 58.01443, 56.88947, 57.08403, 58.79262, 62.98716, 68.70476, 
    73.22769, 74.59242, 73.8849, 73.15436, 73.78822, 74.9845,
  67.95179, 67.00564, 65.72301, 64.93632, 66.17059, 66.82233, 64.64048, 
    63.80264, 62.2719, 61.30988, 58.90459, 59.07368, 64.00903, 70.61009, 
    73.88804, 74.49326, 75.40926, 76.6992, 76.85645, 76.04742,
  90.09764, 90.72139, 91.25752, 91.62565, 92.28006, 92.64742, 92.77328, 
    93.27796, 91.64056, 92.39207, 92.91737, 93.29031, 93.72187, 94.49751, 
    95.00919, 95.13869, 94.56719, 95.01028, 95.32809, 95.502,
  83.85318, 85.33681, 86.87961, 88.5861, 90.21783, 92.04086, 93.59383, 
    94.90946, 92.04279, 92.73958, 93.81758, 94.41714, 95.13055, 95.84274, 
    96.67146, 97.78745, 96.91445, 97.81208, 98.05096, 98.28181,
  85.43948, 87.38397, 89.39732, 91.32227, 92.89687, 94.1954, 95.03278, 
    95.82375, 92.24705, 93.09984, 93.33743, 93.80216, 94.63823, 94.66423, 
    95.29613, 95.60341, 95.39054, 96.27837, 97.16467, 98.16281,
  85.78526, 87.86858, 89.51454, 90.86104, 92.14738, 93.00547, 93.42033, 
    93.90382, 91.7673, 92.65318, 93.68018, 94.90995, 96.15283, 97.6111, 
    98.79482, 99.36933, 99.55042, 99.32982, 98.9877, 97.96564,
  82.02245, 83.77554, 85.47026, 86.49902, 87.64359, 88.32149, 87.89529, 
    87.84527, 86.47792, 86.21529, 86.79842, 88.17248, 90.94182, 93.8168, 
    94.99292, 95.86628, 98.24717, 98.83273, 98.70261, 98.11491,
  82.26412, 83.60612, 84.86308, 85.97424, 87.01152, 87.58945, 87.40823, 
    87.05984, 81.59734, 81.12989, 81.56258, 82.64344, 84.10252, 85.65776, 
    86.82297, 87.86618, 94.48861, 94.88517, 95.07291, 94.53358,
  95.54932, 94.08508, 92.92601, 91.78015, 91.01691, 90.76274, 90.07295, 
    89.71767, 82.08933, 82.37434, 83.47449, 72.23738, 73.53178, 81.07138, 
    86.2747, 81.08817, 87.48873, 89.46902, 90.55835, 91.1777,
  93.83712, 92.63711, 91.02435, 89.89983, 89.50505, 90.20441, 90.98463, 
    91.05991, 84.85093, 85.41405, 88.08123, 84.88241, 85.91866, 90.29426, 
    94.40551, 95.44257, 95.43658, 94.69458, 89.40028, 90.60996,
  68.94599, 69.60528, 70.325, 71.35139, 72.95952, 74.21179, 74.48703, 
    73.17432, 70.51951, 70.04704, 70.74457, 74.91367, 80.06628, 85.0615, 
    86.90202, 88.03505, 91.47592, 93.8731, 96.37093, 95.64284,
  72.06194, 73.60769, 74.2911, 74.13915, 73.75381, 73.36285, 73.6003, 
    74.11332, 75.69495, 76.03605, 76.30199, 76.44465, 76.28757, 75.98466, 
    74.06562, 71.77155, 70.16525, 69.589, 70.03176, 73.74518,
  77.48104, 77.97255, 77.99244, 77.83714, 77.70232, 77.73286, 78.0331, 
    78.37363, 79.27444, 79.71599, 79.75443, 79.79748, 79.69712, 78.77363, 
    76.76929, 74.55019, 72.30096, 70.8222, 70.60889, 71.29136,
  79.31559, 79.80649, 80.35156, 80.94974, 80.81783, 79.47984, 78.94495, 
    80.34335, 82.73627, 83.73847, 83.8989, 83.466, 82.7797, 81.95643, 
    80.25647, 78.37525, 76.4519, 74.45359, 73.06109, 72.86839,
  79.45236, 81.16573, 83.02129, 84.62302, 84.59184, 82.77066, 79.5368, 
    77.5333, 78.26926, 80.14264, 81.26103, 82.09634, 82.94814, 83.54864, 
    84.2702, 84.38338, 83.32738, 81.12894, 78.66229, 76.87337,
  74.85094, 76.90729, 79.94781, 81.46396, 81.00334, 79.38335, 77.48074, 
    76.35844, 76.46294, 77.09204, 77.64252, 79.19589, 81.42252, 83.35685, 
    85.02338, 86.25086, 86.1395, 85.63551, 85.06441, 83.67087,
  70.17616, 71.6972, 74.39901, 76.47809, 77.35523, 77.51985, 77.29112, 
    76.94244, 77.64458, 79.08827, 81.30406, 83.63139, 85.24992, 85.63969, 
    85.14706, 85.09174, 84.27804, 83.62642, 84.40724, 85.2659,
  68.69841, 70.34574, 72.35883, 75.10469, 77.77556, 79.69626, 81.19175, 
    83.01151, 84.58768, 85.3433, 85.93012, 86.28569, 86.2504, 85.57568, 
    83.72828, 82.12981, 80.65338, 79.92384, 81.0628, 81.36863,
  72.95445, 75.7032, 78.89871, 82.08911, 83.98963, 84.85088, 84.91859, 
    84.13863, 82.57323, 82.06425, 82.58173, 83.00074, 83.06938, 82.60606, 
    81.09331, 79.5516, 77.59963, 76.53362, 76.12263, 76.37186,
  80.98055, 83.98367, 87.03001, 87.85546, 86.41217, 83.52869, 80.85545, 
    75.89859, 68.08882, 65.75172, 67.55265, 70.27091, 72.64108, 73.98525, 
    74.86293, 74.85146, 72.8846, 70.25192, 69.15826, 70.17667,
  81.07411, 83.19343, 83.94568, 81.71643, 78.80936, 77.42168, 74.17243, 
    65.39198, 60.65968, 57.78622, 57.06501, 58.31885, 61.12471, 64.67477, 
    68.0128, 69.16209, 68.21843, 67.26512, 68.13016, 70.75298,
  72.83763, 73.30046, 72.85699, 72.02186, 73.00867, 73.4853, 70.75729, 
    71.09572, 69.51138, 66.88995, 61.13041, 59.88748, 63.8336, 67.61614, 
    69.13141, 69.11677, 68.39562, 69.50028, 71.66987, 73.77575,
  91.33452, 91.76824, 92.08362, 92.6461, 93.05537, 93.34305, 93.74966, 
    94.22072, 92.76324, 93.38306, 93.58613, 93.88798, 94.33878, 94.90602, 
    95.38822, 95.11449, 94.72191, 94.8782, 94.91058, 95.01981,
  87.63786, 88.89783, 90.1502, 91.41713, 92.57571, 93.73566, 94.51948, 
    95.18851, 91.76431, 92.50947, 92.71036, 92.91778, 93.13592, 94.369, 
    95.53339, 96.17159, 94.37905, 95.81921, 97.01616, 97.67191,
  89.83316, 91.15501, 92.42437, 93.44006, 94.37505, 95.4507, 95.80059, 
    95.93625, 91.79609, 92.97855, 93.93633, 94.83365, 95.92187, 96.6661, 
    96.92111, 96.40736, 94.99493, 94.91264, 95.77235, 96.53523,
  86.98603, 88.76668, 90.20747, 91.30123, 92.3008, 94.33846, 96.29298, 
    96.97754, 94.63472, 95.2058, 95.71549, 96.06262, 96.3681, 96.62346, 
    96.77101, 97.45914, 97.73247, 97.36315, 96.27975, 95.22832,
  82.83216, 85.03046, 87.52985, 89.66335, 90.95822, 90.99023, 91.6777, 
    92.14835, 92.01165, 93.0901, 94.45315, 95.3533, 96.2709, 96.52122, 
    96.01585, 95.89493, 97.80331, 97.96107, 98.66088, 98.73463,
  83.21659, 85.01691, 85.57825, 85.77547, 86.11076, 86.5942, 86.73833, 
    87.20347, 83.52631, 84.1053, 84.70852, 85.81654, 87.17033, 88.51268, 
    89.23674, 90.29654, 96.71954, 97.78689, 98.03944, 98.14432,
  91.16942, 90.09016, 88.1814, 87.52167, 87.04041, 87.18358, 87.06421, 
    86.94119, 78.82661, 79.55505, 81.7703, 78.53176, 79.64829, 83.32984, 
    85.81514, 83.64087, 88.54162, 90.22079, 91.45371, 91.58527,
  91.14741, 90.72503, 90.58128, 91.11018, 92.07581, 93.67627, 94.74699, 
    95.01267, 89.4548, 89.94464, 91.41414, 86.81541, 86.19673, 88.26128, 
    93.5853, 93.84334, 93.8762, 90.40251, 90.13002, 90.70399,
  78.95053, 78.62708, 83.55924, 88.04285, 88.9893, 89.64762, 90.8205, 
    92.34657, 91.0332, 91.81954, 92.91328, 93.68665, 94.06097, 94.22066, 
    92.89256, 92.51338, 94.70696, 97.07285, 97.01488, 95.55314,
  69.46008, 70.20747, 72.49118, 73.46018, 72.27583, 69.90234, 70.258, 
    71.95185, 73.07703, 73.75069, 75.13992, 75.12772, 74.06981, 72.26141, 
    69.08361, 67.75104, 70.31644, 76.78862, 86.13218, 93.61565,
  71.18409, 73.20511, 74.10941, 73.36915, 71.75227, 70.84105, 70.96215, 
    71.85337, 73.57081, 74.79281, 75.47917, 75.85963, 76.01205, 75.75286, 
    74.6091, 72.90319, 71.73605, 70.39999, 70.19518, 71.6572,
  72.35789, 72.75075, 73.29111, 73.96391, 73.54483, 71.88484, 71.62077, 
    73.31436, 76.51002, 78.8089, 79.99392, 80.55013, 80.51437, 80.13189, 
    79.7942, 78.72033, 77.76295, 76.36597, 74.98575, 74.42455,
  76.10389, 76.6019, 77.08121, 77.40427, 77.48006, 76.30514, 74.08395, 
    72.69298, 74.04079, 76.6266, 78.64362, 80.00111, 81.15939, 82.24097, 
    82.86208, 82.62143, 81.2789, 79.58842, 78.04463, 76.75201,
  73.28427, 73.5237, 74.07048, 74.57598, 74.59143, 74.09592, 73.39168, 
    72.95757, 73.52124, 74.62827, 75.65328, 77.50417, 80.69987, 83.8812, 
    85.72278, 85.74618, 83.94686, 82.45582, 81.56576, 80.59354,
  68.38316, 67.49447, 68.19146, 69.13469, 69.49409, 70.1992, 71.11868, 
    71.95698, 73.6957, 76.44852, 79.52557, 82.66051, 85.89458, 88.05362, 
    88.57645, 88.07819, 86.34194, 84.24113, 83.38407, 83.01408,
  66.26901, 65.83502, 66.16503, 67.38969, 69.20081, 71.84013, 74.50709, 
    77.86394, 83.033, 86.8782, 89.06849, 90.34106, 91.10589, 91.00294, 
    89.55164, 88.12239, 86.55594, 84.52418, 83.83105, 82.46306,
  67.00691, 69.07996, 71.91371, 75.51166, 78.95375, 82.15404, 84.53649, 
    86.10793, 87.1867, 88.53491, 90.06263, 91.15862, 91.66431, 91.19289, 
    89.82567, 88.07773, 85.39725, 82.33486, 79.73489, 77.05778,
  74.7704, 78.68346, 82.79063, 85.81046, 86.68301, 85.6629, 84.08369, 
    79.79738, 73.08722, 71.98983, 74.62851, 78.92401, 82.84008, 84.64065, 
    84.74995, 83.1119, 78.18993, 72.24068, 68.33417, 65.76711,
  78.10748, 80.37218, 82.23807, 81.88117, 79.82626, 78.01415, 73.72053, 
    64.99773, 61.95799, 60.15458, 59.44443, 60.62009, 63.29738, 66.79293, 
    68.83437, 68.59112, 65.81741, 63.33272, 62.91325, 63.77951,
  71.24545, 72.1809, 72.60181, 72.5359, 72.24734, 70.24766, 66.14259, 
    67.04494, 67.18208, 66.05124, 59.90845, 59.0369, 63.712, 67.60802, 
    68.1979, 68.02033, 67.69925, 68.10734, 69.48639, 69.63588,
  91.65794, 92.12198, 92.08334, 92.77003, 93.2541, 93.286, 93.82856, 
    94.26003, 93.09415, 93.8464, 94.25155, 94.64926, 94.9344, 95.33833, 
    95.71553, 95.88094, 95.23533, 95.37359, 95.58719, 95.50046,
  88.3968, 89.70726, 91.01031, 92.39716, 93.50674, 94.60114, 95.57118, 
    96.39342, 93.56018, 94.34951, 94.71899, 95.20913, 96.09931, 96.64265, 
    96.63843, 97.13412, 95.11458, 95.72416, 96.36938, 97.34598,
  90.87503, 92.39645, 93.62802, 94.7043, 95.47087, 96.15776, 96.72097, 
    97.30712, 92.4592, 92.71931, 93.66196, 94.43153, 95.59298, 96.7402, 
    98.09754, 98.58762, 98.41515, 99.12743, 99.27354, 99.36385,
  89.04127, 91.21603, 93.07861, 94.67619, 95.64914, 96.51402, 96.8896, 
    97.36579, 95.50693, 96.91138, 97.58251, 97.68083, 97.7825, 98.13454, 
    99.0172, 99.11309, 99.4229, 99.64176, 99.7985, 99.72855,
  87.68919, 90.74838, 93.17252, 94.94682, 96.01738, 96.96776, 97.82162, 
    98.37659, 98.25336, 98.61408, 98.03719, 96.49596, 95.60352, 96.09229, 
    96.73705, 97.21174, 98.7271, 99.23332, 99.60118, 99.71154,
  86.27883, 89.89754, 92.5754, 94.2609, 95.24816, 95.77198, 95.76675, 
    95.72675, 91.57257, 90.59008, 90.58001, 91.35045, 92.30457, 93.353, 
    94.10517, 94.47997, 97.69482, 97.35623, 97.57537, 98.26995,
  95.03949, 94.0045, 95.13008, 95.96127, 96.02657, 95.85696, 95.85492, 
    95.68275, 88.82127, 87.98329, 87.61988, 83.42518, 85.17785, 90.14491, 
    91.90009, 90.55895, 94.96529, 94.98981, 94.25207, 93.70625,
  96.57985, 97.1338, 97.621, 97.65794, 97.92338, 98.37848, 98.64951, 
    98.58828, 95.25769, 96.05735, 95.43111, 92.10203, 92.08295, 93.31325, 
    95.26558, 95.95519, 96.62885, 96.48474, 93.84599, 93.70355,
  95.19563, 95.78562, 96.1357, 96.47526, 96.95406, 97.25397, 97.547, 
    96.87533, 94.69437, 95.42106, 96.65645, 97.13708, 97.03658, 96.70271, 
    95.66474, 95.63113, 97.04568, 98.461, 98.84753, 98.67113,
  93.39533, 93.46684, 94.22782, 95.40313, 95.59123, 94.31409, 92.02619, 
    91.64915, 93.0064, 93.46439, 93.35876, 92.94624, 91.90657, 88.34534, 
    84.57249, 83.4265, 85.85335, 91.38039, 95.45187, 98.9952,
  94.13924, 94.11552, 94.35142, 94.45163, 89.07214, 80.12948, 75.66328, 
    74.75401, 76.72001, 78.79198, 78.92758, 77.29974, 75.18852, 73.55341, 
    72.60137, 71.61483, 71.21921, 71.12099, 72.32883, 74.89046,
  78.64719, 79.21616, 80.71065, 81.12658, 76.17051, 71.17532, 69.5006, 
    69.91006, 72.21599, 73.86243, 74.83205, 75.52881, 76.15713, 76.92118, 
    77.48337, 77.21686, 76.54132, 75.34051, 73.91902, 72.85513,
  71.14343, 72.93658, 75.00895, 76.23801, 76.29475, 74.5297, 72.11387, 
    70.86074, 72.3191, 74.88904, 76.60111, 77.63366, 78.63711, 80.22759, 
    82.14379, 82.85422, 82.00637, 80.47948, 79.25959, 77.6948,
  68.94957, 69.88037, 71.15166, 72.38249, 72.63554, 72.23999, 71.92322, 
    72.06002, 73.10394, 74.47849, 75.61739, 77.03881, 79.19828, 82.75076, 
    86.66408, 88.42078, 87.69532, 86.5658, 85.48608, 83.9678,
  66.1032, 65.21365, 65.82771, 67.41033, 68.41326, 69.30573, 70.31203, 
    71.08222, 72.84859, 75.00234, 77.35625, 79.98796, 83.18531, 86.93211, 
    89.3259, 89.7857, 88.52094, 86.68999, 85.67384, 84.84765,
  61.97937, 61.11489, 61.19942, 63.30452, 65.78844, 68.3952, 70.9246, 
    73.32544, 77.42642, 81.6974, 85.09613, 87.67405, 89.52384, 90.38952, 
    89.15266, 87.29169, 85.51242, 83.88697, 83.31201, 82.01485,
  60.31191, 60.77276, 62.71341, 67.01497, 71.16327, 74.49552, 77.10242, 
    79.13315, 81.47993, 83.99464, 86.25283, 87.88274, 88.67365, 88.44481, 
    86.78898, 85.08054, 82.75696, 80.26083, 78.20969, 76.05322,
  65.64738, 68.71452, 73.02788, 77.39699, 79.72079, 79.42515, 77.89036, 
    73.14121, 67.48344, 67.45852, 70.49282, 74.67851, 78.10256, 79.92361, 
    80.49801, 79.97781, 75.67896, 70.15986, 66.28669, 64.18756,
  69.97357, 71.96494, 73.99803, 74.3539, 73.53833, 72.69265, 68.49417, 
    60.23383, 59.18622, 59.02003, 59.34024, 60.72142, 63.40349, 66.16481, 
    68.11497, 67.7047, 65.31143, 62.94064, 62.08355, 62.22274,
  65.7878, 66.11272, 66.12112, 65.95279, 66.23715, 65.14915, 61.90971, 
    62.33535, 63.1729, 63.04312, 59.68583, 60.23753, 65.39654, 68.75768, 
    69.491, 69.1801, 68.6109, 68.26974, 68.28575, 68.2654,
  93.70518, 93.98118, 94.2249, 94.5734, 94.99754, 95.2388, 95.50401, 95.7709, 
    94.48863, 95.05081, 95.03638, 95.37113, 95.78835, 95.78324, 95.99773, 
    95.8619, 95.41316, 95.75719, 95.84655, 95.70092,
  85.12473, 86.39916, 87.55338, 88.6837, 89.63049, 90.64378, 91.6398, 
    92.65677, 89.72437, 90.67689, 91.43378, 92.44312, 93.65654, 94.76929, 
    95.69173, 96.5593, 95.86031, 96.59725, 97.37192, 98.00981,
  84.83593, 86.9856, 89.1787, 91.24742, 92.76366, 93.71595, 94.2394, 
    94.82552, 90.63463, 91.44388, 92.31704, 93.49101, 95.25979, 96.57635, 
    97.25601, 98.0061, 97.71506, 98.51454, 99.08251, 99.33304,
  88.76341, 90.76441, 92.45535, 94.07336, 95.23409, 95.90705, 96.5903, 
    97.16705, 95.25014, 96.33564, 97.43206, 98.2342, 98.65756, 99.01987, 
    99.33627, 99.44722, 99.66543, 99.68344, 99.62347, 99.48773,
  86.31908, 89.39733, 91.33521, 92.39639, 93.48109, 94.12691, 94.11551, 
    94.2692, 94.35101, 95.23824, 96.2865, 97.51678, 98.39066, 98.94046, 
    99.14987, 99.13071, 99.99351, 100, 99.91637, 99.73114,
  80.80514, 83.34572, 85.36949, 85.55691, 86.66528, 86.80466, 87.4212, 
    87.99509, 84.36929, 85.38896, 86.81733, 88.51319, 90.47406, 92.27998, 
    93.74374, 94.86552, 98.7457, 99.01744, 99.30259, 99.10144,
  96.28489, 92.03654, 93.11839, 93.38066, 92.39287, 92.19163, 92.17921, 
    91.46821, 82.85644, 81.91869, 82.62421, 78.80415, 80.9087, 88.66699, 
    89.0597, 89.09557, 94.6509, 95.88525, 96.61439, 96.94402,
  99.26674, 98.99717, 99.0393, 98.70087, 98.48048, 98.96253, 99.06977, 
    98.99795, 97.26688, 97.407, 98.10965, 96.93504, 96.79445, 98.51134, 
    98.62493, 99.00657, 97.77195, 97.66165, 92.12209, 93.20724,
  96.91017, 97.50506, 97.7018, 97.45181, 97.5755, 97.87419, 97.75647, 
    97.38259, 95.87627, 96.00642, 96.55659, 97.29914, 98.31058, 98.65697, 
    99.27843, 99.17264, 99.05399, 99.40399, 99.1246, 98.88868,
  94.58678, 95.36331, 96.08253, 96.74921, 96.91602, 96.70319, 96.1405, 
    95.3872, 94.91549, 94.99015, 95.26616, 95.5984, 95.81196, 95.97929, 
    95.57302, 94.37209, 92.62813, 92.1012, 93.77693, 96.23808,
  93.16236, 93.54128, 94.46247, 95.19308, 95.16638, 93.46513, 91.47784, 
    91.05849, 89.92072, 90.56638, 91.16325, 91.11198, 89.8493, 85.59494, 
    77.50992, 68.93499, 60.64864, 56.81988, 56.63053, 60.55947,
  91.27896, 90.80501, 90.60406, 91.06667, 90.40037, 81.67982, 70.57234, 
    66.44256, 68.84846, 71.51748, 71.83332, 71.05956, 71.15198, 71.6463, 
    69.87449, 63.02247, 58.78815, 57.56726, 56.59119, 56.62268,
  70.25851, 70.73203, 71.36246, 72.32716, 72.24174, 67.15667, 60.83553, 
    58.43588, 59.5162, 61.48921, 63.01403, 63.87181, 64.72283, 66.22356, 
    68.76471, 70.06322, 69.90785, 68.8607, 67.58118, 66.33675,
  69.04556, 69.19493, 69.58303, 69.42454, 68.6903, 67.68961, 66.70226, 
    65.99499, 66.32198, 67.41849, 68.38981, 69.50687, 71.04672, 73.42464, 
    77.34251, 79.76242, 79.14723, 78.06803, 77.35647, 76.65428,
  65.79239, 64.7877, 65.28164, 66.10233, 66.13362, 66.13517, 66.33626, 
    66.6995, 67.67908, 69.26882, 71.12657, 73.17137, 75.29264, 77.98986, 
    80.98109, 83.04683, 83.06687, 82.329, 82.26244, 82.58572,
  62.28204, 61.44464, 61.41771, 62.74854, 64.57748, 66.6062, 68.47867, 
    70.2665, 73.46991, 77.32832, 80.23227, 82.15067, 83.77778, 86.06941, 
    86.8483, 86.06485, 84.7865, 83.60629, 83.60693, 83.36036,
  61.67805, 62.51623, 64.36259, 67.37563, 70.32893, 72.59834, 74.67594, 
    76.86958, 79.51675, 82.3327, 84.60355, 86.27304, 87.40363, 88.21258, 
    87.39544, 85.79919, 83.37357, 81.0295, 79.34602, 77.45939,
  66.87434, 70.36089, 74.14293, 77.16069, 78.48688, 78.2634, 77.08985, 
    72.71239, 67.02464, 66.22894, 68.87479, 72.84792, 76.71923, 80.03977, 
    81.66973, 81.35033, 77.89621, 72.4277, 68.64857, 66.32262,
  73.14845, 75.63249, 77.32558, 76.82909, 75.29401, 73.63191, 68.93295, 
    60.82364, 59.42626, 57.84443, 58.47353, 61.11171, 64.43194, 67.75986, 
    70.02013, 69.94599, 67.99144, 66.50624, 66.35001, 66.59253,
  71.63322, 71.76785, 71.04063, 69.76882, 69.51704, 68.182, 64.07148, 
    63.20589, 64.46854, 64.20918, 61.87617, 63.02001, 68.38291, 70.26689, 
    70.72742, 70.70723, 70.79639, 71.55202, 73.13336, 74.16136,
  91.1097, 91.59216, 91.95395, 92.33425, 92.83691, 93.19359, 93.64462, 
    94.28935, 93.00459, 93.67743, 94.12907, 94.55277, 94.91351, 95.12996, 
    95.4977, 95.79382, 95.08646, 95.53324, 95.63914, 96.15374,
  82.87206, 84.34001, 85.94152, 87.51698, 89.10911, 90.62405, 92.03245, 
    93.09047, 90.24945, 91.13017, 91.62518, 92.5163, 93.6971, 94.46577, 
    95.8362, 96.31552, 95.11856, 95.66254, 96.08071, 96.55394,
  84.92297, 86.90975, 88.8327, 90.67767, 92.26612, 93.58691, 94.70672, 
    95.46197, 91.281, 92.69986, 94.13078, 95.35294, 96.37712, 97.21168, 
    97.71515, 98.17539, 97.52463, 97.87846, 98.05789, 98.24858,
  87.17742, 89.24651, 91.15928, 93.30486, 94.79043, 95.94138, 96.72774, 
    97.60007, 95.90729, 96.81484, 97.76214, 98.37276, 98.62583, 98.64053, 
    98.65599, 98.61399, 98.73685, 98.74942, 98.90218, 99.17446,
  84.08456, 86.3009, 88.04773, 89.61918, 91.07851, 92.32195, 92.76308, 
    93.22322, 93.05325, 94.25188, 95.26844, 96.77962, 97.94419, 97.96227, 
    97.69012, 97.34319, 98.30791, 98.56308, 98.84583, 98.53413,
  82.80671, 84.78013, 86.38032, 87.69786, 87.97816, 88.30051, 88.06248, 
    88.6033, 84.63933, 85.51894, 86.88718, 88.41724, 90.08943, 91.19088, 
    91.73224, 92.07465, 96.95744, 98.17738, 98.85744, 98.36217,
  95.23962, 94.76284, 94.78583, 94.47859, 93.23164, 92.05632, 90.89611, 
    90.46159, 82.60683, 82.80305, 84.12147, 77.88493, 79.26337, 85.53088, 
    87.0089, 85.18975, 91.66454, 94.12804, 95.18323, 95.03426,
  97.73817, 97.67179, 97.75729, 97.72355, 97.33146, 96.53381, 95.82396, 
    95.94714, 92.87679, 93.74361, 94.52656, 92.47122, 92.32223, 94.21955, 
    96.38732, 97.70341, 96.5364, 93.81056, 89.85317, 90.29899,
  97.9027, 98.03225, 98.38633, 98.68135, 98.76539, 98.53503, 98.37715, 
    97.91383, 95.15115, 95.20081, 95.78004, 96.50418, 97.12886, 97.14656, 
    97.27493, 97.64686, 98.3799, 98.93739, 98.42317, 98.58811,
  97.28354, 97.28559, 97.56422, 97.63713, 97.62814, 97.65409, 97.08708, 
    96.16943, 95.5517, 95.28419, 95.83575, 95.83221, 95.82552, 95.74289, 
    95.84385, 96.19891, 95.38385, 94.8995, 94.18235, 94.36251,
  96.17837, 96.2021, 96.21857, 96.08974, 96.06056, 95.75645, 95.41219, 
    94.66755, 94.5983, 94.92978, 95.46617, 95.80333, 95.78063, 95.30835, 
    94.88222, 94.27081, 90.21914, 83.06027, 76.71523, 75.92358,
  92.89462, 92.05207, 91.59364, 91.66467, 92.72347, 91.73662, 88.55994, 
    85.23506, 85.20387, 87.44485, 90.08914, 90.50726, 90.29597, 90.67332, 
    92.01646, 91.31819, 84.73391, 75.69726, 66.15163, 62.22515,
  77.70807, 78.45634, 79.86636, 81.52048, 83.04637, 82.37428, 78.80828, 
    75.25638, 75.04809, 76.60947, 77.99258, 78.44479, 78.33889, 78.16547, 
    79.43428, 80.11105, 77.06127, 72.60514, 68.76777, 66.62313,
  73.23197, 74.74776, 76.13705, 76.99931, 77.07592, 76.41173, 75.24165, 
    74.21696, 74.1329, 75.54197, 76.71712, 77.72709, 78.53407, 79.08987, 
    80.4119, 81.45206, 79.21304, 76.98203, 75.44963, 74.04202,
  70.56814, 70.28458, 70.67419, 71.24238, 71.25203, 71.40958, 71.57849, 
    71.87988, 72.62862, 74.47387, 76.6801, 78.77718, 80.2541, 81.18396, 
    82.21152, 83.44368, 82.86115, 81.24197, 79.85084, 79.35873,
  67.62677, 67.05627, 66.66162, 67.46214, 69.04508, 71.14854, 72.91283, 
    74.3063, 76.18599, 78.9655, 81.29922, 82.5677, 83.62609, 85.53981, 
    87.38722, 87.18274, 85.028, 82.75948, 81.41428, 79.72343,
  65.8767, 66.87949, 69.00241, 72.08866, 74.85966, 76.95855, 78.60165, 
    80.2327, 81.59835, 83.342, 84.68747, 85.45665, 86.07793, 87.01159, 
    87.13952, 85.43329, 81.87719, 78.35767, 75.60091, 72.75599,
  71.89007, 75.65775, 79.49545, 82.33424, 83.25751, 83.10851, 82.47941, 
    78.42627, 73.28499, 72.07269, 72.81808, 74.44689, 76.55704, 78.58655, 
    79.2086, 77.96556, 73.31664, 67.75738, 63.64846, 61.05314,
  81.35389, 84.4427, 85.82452, 84.99022, 83.43957, 83.23944, 80.64889, 
    72.85186, 70.37888, 67.17081, 65.18749, 65.26502, 66.07677, 66.31205, 
    66.16408, 65.09998, 62.22377, 59.8134, 58.83548, 59.09148,
  82.51872, 82.98526, 81.65105, 79.75537, 79.79219, 79.63465, 74.36787, 
    67.25586, 69.31104, 68.9579, 66.78568, 66.27446, 69.73946, 68.99075, 
    66.43671, 65.18057, 64.74754, 65.02265, 66.41135, 68.00977,
  92.53941, 92.92354, 93.42612, 93.50632, 93.8541, 94.29669, 94.56229, 
    94.68472, 93.16457, 93.55772, 93.75191, 93.9202, 94.2494, 94.49371, 
    95.01101, 95.05447, 94.26254, 94.60038, 94.80488, 95.04651,
  86.46848, 87.40259, 88.49599, 89.61371, 90.70206, 91.79354, 92.81082, 
    93.77392, 90.36663, 91.62245, 92.53781, 93.48852, 94.35068, 95.31064, 
    96.29751, 97.02515, 95.31661, 95.95338, 96.5107, 97.0204,
  84.46863, 86.01861, 87.50409, 89.22029, 90.64022, 92.11431, 93.36309, 
    94.73772, 90.57343, 91.62907, 92.65103, 93.3326, 94.20158, 95.17296, 
    95.95168, 96.49588, 94.87959, 95.62034, 96.37105, 96.83612,
  84.52866, 86.58179, 88.13055, 89.8911, 91.6841, 93.27789, 94.94929, 
    96.4386, 94.7424, 95.75379, 96.53352, 97.06603, 97.35815, 97.52422, 
    97.60863, 97.4486, 97.894, 98.07104, 98.05618, 97.89325,
  81.58457, 83.51334, 85.29884, 86.91253, 88.45502, 90.01276, 91.39989, 
    92.74631, 92.36508, 94.05685, 95.01661, 95.31708, 95.81408, 96.34525, 
    96.40888, 96.28043, 98.8241, 98.66712, 98.24263, 97.32677,
  82.37822, 84.35499, 86.13895, 87.24657, 87.74308, 88.15745, 88.16116, 
    87.78851, 83.9006, 84.40176, 85.09687, 86.13441, 87.43996, 88.77401, 
    89.93854, 91.19897, 97.31217, 97.6596, 97.76043, 97.34863,
  92.35216, 90.98985, 90.95733, 91.49788, 92.04906, 92.11428, 91.89627, 
    91.51053, 83.40427, 83.45, 84.22855, 78.62718, 79.10769, 84.51613, 
    87.24924, 85.43359, 92.1765, 94.34116, 95.61265, 95.7862,
  95.05501, 94.2516, 92.92873, 93.44405, 94.535, 94.77725, 95.40251, 95.307, 
    91.35632, 92.0526, 92.66164, 89.59322, 89.93682, 93.40008, 96.34988, 
    96.17606, 96.77372, 95.02788, 94.2688, 95.54061,
  97.46338, 97.2522, 96.80891, 96.28575, 95.72438, 95.25581, 94.98406, 
    94.85722, 93.07681, 93.63505, 94.13689, 94.32594, 94.23279, 94.41785, 
    94.76115, 95.28768, 95.97369, 96.5938, 96.06327, 96.54994,
  95.73717, 95.87534, 95.89588, 96.05107, 95.92085, 95.73313, 95.32261, 
    95.00114, 94.79707, 94.79238, 94.62641, 94.36758, 94.16814, 94.03672, 
    94.62723, 95.68829, 96.29477, 96.78045, 96.54723, 95.99476,
  94.73631, 94.61339, 94.40717, 94.10931, 94.14356, 94.00336, 93.63068, 
    93.2951, 92.67144, 92.58344, 92.59695, 92.66691, 92.69752, 92.80316, 
    92.98133, 93.14464, 93.13647, 93.0798, 92.38663, 90.57652,
  94.14833, 93.46005, 92.43086, 91.87246, 91.77451, 91.40665, 89.81047, 
    86.86695, 84.29136, 83.28316, 82.76315, 82.38354, 82.12502, 83.29446, 
    85.28006, 86.08701, 86.13319, 84.98151, 80.86469, 75.50568,
  87.59497, 86.74735, 86.07873, 84.81692, 83.45614, 81.17982, 76.63614, 
    71.76033, 70.59795, 71.8457, 72.83611, 73.54501, 74.17467, 75.17702, 
    77.39095, 79.26134, 79.38712, 77.90476, 75.52119, 73.51862,
  79.19885, 79.45852, 79.48485, 78.39234, 76.54414, 74.1515, 71.9894, 
    70.6656, 70.4724, 71.51627, 72.77909, 74.31207, 76.08923, 78.33427, 
    81.14893, 83.25776, 82.73442, 81.86871, 81.09628, 79.95679,
  75.67793, 73.74133, 73.21755, 72.95041, 72.01845, 71.12457, 70.57544, 
    70.22608, 70.35497, 71.5131, 73.39555, 75.9522, 78.36761, 80.21629, 
    81.61873, 83.21422, 84.11247, 84.12509, 84.10716, 84.71982,
  70.65956, 68.64211, 67.4321, 67.18739, 67.85838, 69.43364, 71.133, 
    72.45114, 74.11443, 76.44806, 78.90216, 81.14935, 83.05303, 84.86434, 
    86.31036, 86.73701, 86.13105, 85.13618, 85.27533, 84.9712,
  67.69324, 67.06417, 67.41206, 69.12985, 71.30246, 73.41824, 75.44501, 
    77.12562, 78.75966, 80.86021, 83.09206, 84.44192, 85.17146, 86.01516, 
    85.99961, 85.10615, 83.16496, 81.18698, 79.52399, 77.50517,
  69.29246, 71.38155, 74.40289, 76.95641, 77.96749, 77.76231, 77.18858, 
    72.39681, 66.53722, 65.17691, 67.35666, 71.53838, 74.94732, 77.09969, 
    77.97482, 77.46228, 74.76048, 70.59315, 67.95928, 67.02927,
  72.55556, 74.31676, 75.79509, 74.85108, 72.93807, 71.35282, 67.43378, 
    60.07803, 55.88239, 54.0007, 54.90176, 57.38945, 60.51659, 63.30316, 
    66.43961, 68.17341, 67.54629, 66.84351, 67.52925, 68.96636,
  69.26862, 69.01531, 67.89384, 65.95235, 64.82139, 63.73297, 61.11056, 
    62.39193, 64.2748, 64.05579, 60.35431, 58.71916, 62.88017, 65.91654, 
    69.25653, 71.80682, 73.53966, 74.74963, 76.36543, 77.74026,
  91.53083, 91.86279, 92.15949, 92.39041, 92.63016, 92.90179, 93.16399, 
    93.48732, 91.9562, 92.2211, 92.43272, 92.66709, 92.96333, 93.2302, 
    93.44633, 93.61163, 92.74581, 92.872, 93.16305, 93.33115,
  86.3987, 87.17014, 88.01995, 88.77533, 89.82421, 90.61562, 91.45008, 
    92.46239, 88.80419, 89.63085, 90.26646, 90.92902, 91.58669, 92.32581, 
    93.11859, 93.89718, 91.90701, 92.58995, 93.21559, 93.71144,
  83.74517, 85.00637, 86.18618, 87.40044, 88.57651, 89.69822, 90.90589, 
    92.09085, 87.69324, 88.82745, 89.92931, 90.7478, 91.78677, 92.769, 
    93.66597, 94.54227, 92.29524, 93.43977, 94.1682, 94.75268,
  84.72129, 86.09185, 86.92377, 87.48589, 88.78668, 90.31037, 91.58701, 
    92.89511, 90.58941, 91.52543, 92.8584, 93.94341, 94.77242, 95.38774, 
    95.90946, 95.93398, 96.49706, 96.40445, 96.27139, 96.1813,
  83.56911, 85.12084, 86.57307, 86.67006, 87.66581, 88.89671, 89.99959, 
    90.63262, 89.4394, 90.17187, 91.22892, 92.15958, 93.29126, 94.2504, 
    94.73612, 94.68822, 98.3769, 98.2146, 97.8203, 97.0973,
  81.93482, 84.13534, 85.16996, 85.8568, 86.3764, 86.21828, 85.66315, 
    85.59066, 81.20061, 81.76836, 82.3584, 83.68143, 85.25578, 87.08389, 
    88.96532, 90.77719, 97.63326, 98.06855, 98.0603, 97.51938,
  89.20885, 87.02596, 86.56017, 86.64511, 86.48782, 86.04251, 85.44414, 
    84.89719, 76.67503, 76.36691, 75.58459, 73.57614, 75.37121, 81.59487, 
    84.00529, 83.8856, 91.87019, 94.74844, 96.36301, 96.98526,
  94.82829, 93.13435, 92.10718, 91.60255, 91.39457, 91.45196, 91.6768, 
    91.76466, 87.7364, 87.00246, 84.09727, 85.63181, 86.59966, 91.03868, 
    91.87273, 88.93357, 89.63835, 91.92227, 90.43349, 92.94894,
  96.00591, 95.86395, 95.52243, 94.75134, 94.01276, 93.73091, 93.40109, 
    92.84409, 90.93029, 90.88951, 90.43187, 89.23586, 89.36074, 90.29819, 
    91.63103, 91.95956, 90.09693, 91.42274, 91.52522, 93.20019,
  95.51899, 95.17882, 95.41393, 95.34388, 95.29506, 95.11456, 94.8427, 
    94.10665, 93.3046, 92.73495, 92.24863, 91.56606, 91.05747, 91.22786, 
    91.95469, 93.02588, 93.46126, 93.36666, 93.72321, 93.96754,
  96.50563, 95.98273, 95.72543, 95.647, 95.50613, 95.3802, 95.31524, 
    94.91688, 94.04503, 93.53355, 93.0673, 92.74772, 92.45072, 92.516, 
    92.42985, 92.10853, 91.72982, 91.74052, 91.64668, 91.48965,
  95.40668, 95.5597, 95.74107, 95.85821, 95.82025, 95.52161, 94.94604, 
    94.18866, 92.6305, 91.98547, 91.45533, 90.81157, 90.15099, 89.85983, 
    89.78664, 89.37697, 87.68431, 85.56686, 76.78193, 68.49215,
  92.41322, 92.9977, 93.08356, 92.52613, 91.64633, 89.70079, 85.76343, 
    82.00089, 79.74434, 79.1631, 78.2567, 77.21842, 75.99715, 74.73933, 
    74.07844, 73.80713, 71.04377, 67.29123, 64.30585, 63.30486,
  87.4014, 88.3419, 89.01124, 88.84686, 87.22945, 84.79037, 81.96977, 
    79.84908, 77.8607, 77.46011, 76.7327, 76.2067, 75.78065, 76.07384, 
    76.7852, 76.84704, 73.6523, 71.80834, 71.60554, 71.57381,
  82.26418, 82.01357, 82.74786, 83.68079, 83.32159, 82.36074, 80.72399, 
    78.61414, 75.96603, 75.52299, 75.95756, 76.87415, 77.33549, 77.48283, 
    77.31706, 76.98409, 75.49948, 75.2066, 76.12678, 77.74934,
  77.03176, 76.80267, 77.17622, 77.9864, 78.36169, 78.43922, 78.01104, 
    76.8017, 75.2916, 76.00603, 77.19794, 77.69083, 77.76075, 78.10917, 
    79.13309, 79.5898, 78.04587, 76.64787, 76.85881, 76.78043,
  74.16988, 75.26602, 75.51107, 75.41006, 75.0127, 74.84903, 74.55793, 
    74.69054, 74.76961, 75.75549, 76.50631, 76.62746, 76.49383, 76.8923, 
    77.73635, 77.77654, 75.06453, 72.29245, 70.3081, 68.49146,
  75.01647, 76.52116, 76.99572, 75.93379, 74.09873, 72.94416, 72.89487, 
    70.7845, 66.86546, 65.88825, 66.41423, 67.43385, 68.74383, 70.04481, 
    71.21117, 71.09162, 67.57551, 63.85808, 62.11641, 61.98838,
  75.80585, 75.00981, 72.16908, 70.76083, 70.95772, 73.08678, 72.41461, 
    67.57222, 63.25515, 59.67884, 57.70361, 57.46632, 58.60918, 60.16326, 
    61.1398, 60.46657, 58.6221, 58.51988, 59.90939, 61.88026,
  70.29688, 68.10478, 65.51565, 66.70145, 70.19799, 72.85743, 71.65115, 
    70.37383, 70.65482, 68.18252, 63.56903, 60.03951, 62.25284, 64.39246, 
    64.18719, 63.62231, 62.49077, 62.73181, 64.22783, 65.69978,
  93.40524, 93.63052, 93.74477, 93.92133, 94.07227, 94.36821, 94.56038, 
    94.79021, 93.15051, 93.3344, 93.53109, 93.6391, 93.75005, 93.91359, 
    94.17525, 94.25866, 93.1165, 93.35694, 93.3438, 93.47266,
  87.34984, 87.93036, 88.55212, 89.24193, 89.7633, 90.49643, 91.33537, 
    92.34826, 88.81252, 89.7149, 90.51307, 91.27046, 91.86879, 92.36327, 
    92.63201, 93.56127, 91.55492, 92.06484, 92.25854, 92.67072,
  83.01681, 84.65521, 85.83791, 86.69213, 87.65654, 88.79309, 90.01127, 
    91.11053, 86.97298, 87.76248, 89.12636, 90.49484, 91.29797, 91.9342, 
    92.44392, 93.3428, 91.09727, 90.89201, 91.21043, 91.23952,
  83.01707, 84.71975, 86.33137, 87.78274, 88.86682, 89.86069, 90.75421, 
    91.81506, 89.2961, 89.84932, 90.6769, 91.57087, 91.75528, 92.03206, 
    92.44347, 92.66174, 93.33704, 93.13696, 92.7206, 92.08897,
  82.74805, 85.13705, 87.04423, 88.58694, 90.39852, 91.58619, 92.5016, 
    93.08026, 91.78036, 92.45865, 92.79546, 92.84111, 93.60711, 93.73257, 
    93.70904, 93.46683, 97.54133, 97.44352, 97.45401, 97.25115,
  82.19572, 84.83828, 86.86433, 88.22082, 89.2732, 90.07162, 90.8071, 
    91.37184, 87.41505, 87.64985, 88.0142, 88.49524, 89.10714, 89.85517, 
    90.79215, 91.84208, 98.06209, 98.30605, 98.69833, 98.43236,
  88.23204, 86.40644, 85.95792, 86.45122, 86.46683, 86.11591, 85.55882, 
    84.85355, 76.88212, 76.00072, 74.86147, 76.83327, 78.5031, 82.2042, 
    84.34595, 86.6403, 94.20827, 96.06183, 97.11873, 97.24681,
  92.93485, 93.31217, 93.74967, 93.84625, 93.56619, 92.9314, 92.13322, 
    91.38534, 83.99986, 81.47729, 77.66013, 81.40992, 82.26608, 86.81381, 
    81.9156, 77.55446, 79.83798, 92.241, 92.26324, 93.92339,
  93.64618, 92.88976, 92.64704, 92.45972, 92.34485, 92.27419, 92.28371, 
    92.44556, 90.05258, 89.61297, 88.97463, 89.02045, 89.54876, 89.7478, 
    90.97975, 92.01121, 92.16415, 90.90589, 93.01569, 94.9967,
  95.71848, 94.76565, 93.62211, 93.41756, 93.75989, 94.48754, 95.34542, 
    95.52589, 95.07485, 94.55515, 94.7486, 95.64413, 96.18783, 96.30763, 
    96.16676, 96.1309, 96.37945, 96.6591, 96.97069, 97.03493,
  93.90414, 93.51788, 92.95254, 92.05329, 91.77734, 92.26482, 92.9285, 
    93.2967, 93.48712, 93.36066, 93.20174, 93.57171, 94.46699, 94.89774, 
    94.40071, 93.56737, 93.73723, 94.20942, 94.50231, 94.53419,
  88.81693, 88.37515, 88.01591, 88.30602, 88.562, 88.70956, 88.6641, 
    88.97151, 89.4008, 89.21641, 88.86186, 89.28584, 90.3072, 91.34736, 
    91.86616, 90.83864, 90.92561, 90.93531, 90.00346, 89.19898,
  89.43542, 89.13025, 88.49283, 88.04377, 88.05888, 87.54561, 85.24924, 
    83.21009, 82.98197, 83.71181, 83.99631, 84.58853, 85.68697, 87.08511, 
    89.06136, 90.58186, 91.89162, 91.71532, 91.11156, 89.70659,
  84.47961, 84.68265, 84.92085, 84.35423, 83.10053, 81.68184, 80.00011, 
    78.50604, 77.83684, 78.46842, 79.61284, 81.09853, 82.86624, 85.24609, 
    88.72567, 91.45831, 92.45761, 92.75439, 93.6637, 93.42393,
  78.72286, 77.18143, 76.88543, 76.7821, 76.17042, 75.58565, 75.10949, 
    74.89845, 75.64461, 77.36304, 79.32475, 81.69822, 84.11619, 86.36036, 
    88.56317, 89.7836, 90.43902, 91.1668, 92.80505, 93.97121,
  75.44806, 73.93626, 73.05721, 73.22399, 73.73972, 74.61746, 75.65232, 
    77.00131, 78.5237, 80.56525, 82.81727, 84.61097, 86.25597, 87.88342, 
    88.94178, 89.31367, 89.39072, 89.26147, 90.64751, 91.45557,
  74.55026, 74.60702, 75.05669, 75.79292, 76.80929, 77.59938, 78.31848, 
    79.05762, 79.49974, 80.50008, 82.00977, 83.2114, 84.52235, 86.10838, 
    86.84188, 87.14774, 86.07437, 84.99219, 85.0402, 84.62097,
  77.02428, 77.92416, 78.42152, 78.53931, 78.42303, 78.04944, 77.24231, 
    73.36998, 68.25177, 67.71845, 69.52915, 72.98062, 76.18314, 78.70367, 
    80.296, 80.73996, 78.91735, 76.03487, 74.29453, 73.13023,
  80.69221, 80.64408, 78.94405, 76.3064, 74.08175, 72.66514, 68.86243, 
    63.33049, 59.16113, 56.28193, 56.26172, 59.21124, 64.06935, 67.17268, 
    69.35572, 70.06043, 68.62807, 67.03411, 67.53008, 69.8196,
  76.51835, 75.86806, 73.67548, 70.73037, 69.21645, 67.47099, 64.106, 
    61.12835, 60.23363, 59.21764, 59.35999, 60.45935, 66.60027, 70.1373, 
    70.02644, 69.25018, 68.09383, 68.62275, 71.62584, 75.71154,
  92.44301, 92.55415, 92.81008, 93.07385, 93.29446, 93.47301, 93.57725, 
    93.81602, 92.35689, 92.40112, 92.55384, 92.80453, 92.9448, 93.13641, 
    93.19223, 93.38131, 92.68352, 92.89144, 93.01014, 93.1354,
  85.90691, 86.56623, 87.23544, 87.94296, 88.85885, 89.74689, 90.85666, 
    91.75288, 88.25063, 88.74602, 89.43264, 90.28096, 90.82127, 91.33741, 
    91.96165, 92.46669, 90.32439, 90.62839, 91.21921, 91.56152,
  83.38426, 84.42619, 85.23798, 86.00578, 86.86459, 87.85238, 88.84778, 
    89.92807, 85.67677, 86.73628, 87.56963, 88.73261, 89.65799, 90.48551, 
    91.01672, 91.54141, 89.59077, 90.17033, 90.55505, 91.10084,
  83.9388, 85.16045, 86.01005, 86.83165, 87.52094, 88.30606, 89.28807, 
    89.66106, 86.38295, 87.17905, 88.4113, 89.17462, 89.63024, 90.31876, 
    90.77094, 91.05009, 92.02879, 92.83823, 93.35644, 93.28868,
  83.7319, 85.45763, 86.74174, 87.90202, 89.35737, 90.73767, 91.88318, 
    92.26033, 90.74712, 90.65824, 91.01485, 90.96249, 91.14425, 91.18721, 
    91.2074, 91.39996, 95.68079, 95.61222, 95.70278, 95.39819,
  83.4076, 85.727, 87.85223, 89.37799, 90.63172, 91.21497, 91.54541, 
    91.76778, 87.81484, 87.63295, 88.01273, 88.40845, 89.24387, 90.2965, 
    91.3476, 92.05641, 97.936, 97.66911, 97.19583, 96.57883,
  89.16943, 86.72224, 85.92068, 86.42038, 86.23916, 85.73095, 85.152, 
    84.45525, 75.93121, 74.86727, 74.40192, 76.3188, 78.16763, 82.61976, 
    83.28049, 85.75433, 92.92856, 94.80295, 95.66848, 95.89293,
  91.89663, 91.30896, 89.68515, 86.3188, 83.1523, 80.30015, 78.34389, 
    76.22459, 68.21365, 66.71136, 66.94849, 72.87475, 73.4457, 75.05812, 
    65.92447, 69.72328, 74.82589, 91.1685, 92.29793, 93.88995,
  86.99989, 86.91304, 87.02068, 86.43614, 85.04331, 83.59402, 81.66628, 
    79.37112, 75.37344, 74.2392, 74.36598, 75.28647, 77.78413, 81.52263, 
    85.88183, 88.58099, 88.49821, 86.22623, 90.47041, 93.95533,
  88.88998, 88.41317, 88.29765, 87.35829, 86.19786, 85.03641, 83.86858, 
    82.46651, 80.94958, 80.3077, 81.15719, 82.32502, 82.89332, 83.8418, 
    85.83334, 88.82185, 90.92731, 92.31435, 93.24147, 93.95045,
  87.15033, 87.84296, 87.72257, 86.76282, 85.60578, 85.07864, 85.14627, 
    85.83188, 85.66997, 83.96107, 83.09772, 83.32456, 83.81047, 83.45884, 
    82.8449, 83.39531, 84.38712, 85.73657, 86.81988, 88.31633,
  86.7394, 86.70347, 87.21224, 87.83609, 87.99838, 87.23609, 86.41866, 
    86.97437, 88.79739, 88.20078, 86.08281, 84.39985, 84.07814, 84.48129, 
    84.93804, 85.30326, 85.67323, 85.97694, 85.43481, 85.24931,
  88.26688, 89.00607, 89.58652, 89.53969, 88.55025, 86.26707, 83.21397, 
    82.29993, 83.33906, 84.76199, 84.79298, 83.54269, 83.0423, 84.21339, 
    86.13208, 87.97232, 88.17857, 87.8054, 87.25203, 86.021,
  83.74461, 83.8362, 84.46854, 84.22622, 82.17733, 79.4481, 77.5826, 
    77.23801, 77.80474, 79.1656, 80.64503, 81.6907, 82.82734, 84.35868, 
    86.69841, 88.60161, 88.97796, 89.15794, 89.88519, 90.01824,
  81.5277, 79.20546, 78.33659, 77.89895, 76.764, 76.07089, 75.93476, 
    76.07051, 76.55405, 78.50878, 81.03346, 83.39197, 85.97395, 87.65118, 
    88.35034, 88.87852, 88.9731, 88.59158, 89.94469, 91.49586,
  81.03574, 79.1441, 77.80096, 77.43678, 77.41637, 78.34676, 79.39043, 
    80.11768, 80.74838, 82.33295, 84.2513, 86.10355, 88.15987, 89.62315, 
    89.51392, 88.8745, 88.1041, 87.0652, 88.0163, 88.9641,
  80.7386, 80.66492, 80.73909, 81.17932, 81.36298, 81.74024, 82.106, 
    82.25259, 82.25548, 82.77183, 83.80997, 84.94102, 86.10986, 87.365, 
    87.57264, 86.9896, 85.62181, 83.60249, 82.56335, 82.39453,
  80.87868, 81.95775, 82.87517, 82.40625, 81.47968, 80.72807, 79.88604, 
    76.47758, 71.60101, 70.5452, 72.60847, 75.91441, 78.67392, 80.32207, 
    81.41126, 81.33678, 79.06622, 76.31175, 75.21376, 75.818,
  78.56929, 78.79191, 77.94722, 76.3688, 75.1636, 74.17882, 70.88177, 
    65.40033, 61.60563, 59.56934, 59.96348, 62.39433, 66.21, 69.89199, 
    72.21029, 72.8725, 72.12387, 71.78223, 73.15955, 75.18934,
  69.18991, 68.95726, 68.14276, 68.06258, 69.27203, 68.78416, 65.73855, 
    62.31605, 62.01057, 62.35017, 63.22859, 64.30751, 69.19249, 72.71992, 
    73.53517, 72.98431, 72.48734, 72.99763, 74.73824, 75.69361,
  91.325, 91.62498, 91.91856, 92.11496, 92.36486, 92.6489, 93.03619, 
    93.22375, 91.79601, 92.23297, 92.21837, 92.71189, 92.95911, 93.39848, 
    93.6113, 93.80059, 92.96815, 93.118, 93.25391, 93.27822,
  85.65299, 86.71307, 87.85952, 88.98536, 89.97103, 91.07632, 92.08691, 
    92.90121, 89.49309, 90.55045, 91.38802, 92.19384, 92.86543, 93.53723, 
    94.3108, 95.19808, 93.24117, 94.10963, 94.66381, 95.07856,
  84.52646, 85.73663, 86.90998, 88.24065, 89.66509, 91.12228, 92.77014, 
    94.23345, 90.26763, 91.92609, 93.38231, 94.71088, 95.33937, 95.83434, 
    96.46557, 97.13651, 95.7272, 96.35423, 96.8961, 97.21428,
  83.79275, 85.49293, 87.10849, 89.00546, 90.91644, 92.55302, 93.81554, 
    94.97108, 93.10599, 94.16704, 95.06294, 95.80434, 96.12996, 96.65532, 
    97.14828, 97.57996, 98.54806, 98.51258, 98.35493, 98.15579,
  82.176, 84.51993, 87.00098, 88.94467, 91.10825, 92.70121, 93.61533, 
    94.07767, 92.99275, 93.66022, 94.23866, 94.72334, 95.06922, 95.51804, 
    95.83141, 95.82664, 98.36261, 98.27786, 97.89091, 97.2163,
  80.96848, 83.1399, 84.85093, 86.707, 88.07519, 88.88721, 89.18014, 
    88.96542, 84.71703, 85.40695, 85.83326, 86.93398, 88.06453, 89.4586, 
    90.74474, 91.82777, 97.46333, 97.58763, 97.52428, 97.27587,
  86.42242, 84.56783, 83.6535, 83.69064, 83.63763, 83.85336, 83.90754, 
    83.77508, 76.14974, 75.6136, 74.36138, 74.24282, 76.46488, 83.24268, 
    86.96643, 84.67218, 91.8949, 93.9471, 95.16621, 95.79187,
  82.0963, 78.79285, 75.8448, 73.03033, 71.13911, 70.17095, 69.38113, 
    68.28526, 61.57974, 58.8863, 57.80584, 68.24312, 75.69369, 84.93351, 
    82.60912, 83.67823, 88.31241, 92.52781, 92.36469, 93.35764,
  82.09239, 81.83034, 82.80064, 84.08085, 84.27807, 84.46941, 84.29327, 
    83.77042, 81.10189, 80.83086, 80.40411, 80.09741, 82.172, 85.16044, 
    87.49454, 87.77973, 86.57967, 83.99455, 89.27711, 92.46007,
  88.11375, 87.93916, 88.11992, 88.41995, 88.36337, 88.37748, 88.92747, 
    89.4249, 89.7613, 89.70148, 89.61591, 88.93709, 87.86115, 86.75962, 
    86.04221, 86.4631, 87.38915, 88.93379, 90.20241, 90.77029,
  90.3673, 89.83743, 89.74417, 89.48362, 89.16594, 89.31287, 90.14939, 
    91.08649, 92.04797, 91.92516, 91.57193, 91.166, 90.74265, 89.77627, 
    88.68081, 88.11619, 88.26632, 88.85135, 89.18601, 89.73842,
  88.18355, 87.95055, 88.29538, 88.6764, 88.33576, 87.40854, 87.65707, 
    89.53069, 92.09475, 92.91373, 92.02163, 90.66851, 90.10159, 90.26154, 
    90.14081, 90.07284, 89.71739, 89.14067, 88.12697, 87.14636,
  87.13589, 88.15541, 88.99352, 89.3412, 88.75476, 86.8118, 84.6143, 
    84.35153, 86.56256, 88.44894, 89.21167, 89.25611, 89.05747, 89.37659, 
    90.45618, 91.37931, 90.44997, 89.19081, 88.25457, 86.0503,
  84.52124, 85.01393, 85.92559, 86.35941, 85.70811, 84.36646, 83.22486, 
    82.95805, 83.64801, 84.4488, 85.1534, 86.43736, 87.4975, 88.44962, 
    89.65621, 90.19811, 88.88039, 88.16209, 87.9463, 86.75463,
  81.84708, 80.11159, 80.01262, 80.56998, 80.74506, 81.10082, 82.22531, 
    83.60764, 84.98487, 85.88754, 86.62501, 87.80793, 88.97485, 89.80492, 
    89.80434, 89.32128, 87.93919, 87.0434, 87.40618, 87.88209,
  77.47684, 76.54875, 76.77071, 78.45528, 80.39217, 82.37766, 84.43672, 
    86.17806, 87.66307, 88.73548, 89.4807, 90.36632, 91.3638, 91.27776, 
    90.19287, 89.34803, 87.99957, 87.16957, 87.47681, 87.1743,
  73.99126, 75.50745, 77.76992, 80.43286, 82.49008, 83.8263, 84.36548, 
    85.33559, 86.97656, 87.92945, 88.47642, 88.856, 89.4482, 89.2869, 
    88.80557, 88.2409, 86.43758, 85.04674, 84.10149, 82.97558,
  75.7392, 78.01038, 80.9461, 82.01971, 81.71661, 81.46439, 81.08431, 
    79.68206, 77.92877, 77.74698, 79.40424, 81.76195, 83.72998, 84.80029, 
    84.98946, 84.40895, 82.04494, 79.69085, 78.3793, 77.78555,
  77.12815, 77.75439, 77.19624, 76.36654, 76.51052, 77.04877, 74.60466, 
    70.7486, 67.9005, 65.49918, 65.67699, 68.26649, 71.92208, 75.00044, 
    76.25137, 75.9989, 74.84174, 73.46321, 73.07743, 72.25179,
  71.23436, 69.80621, 67.92341, 68.85827, 71.7654, 72.47925, 70.29117, 
    65.18519, 64.00188, 63.78293, 63.66858, 64.47598, 69.40471, 73.21999, 
    73.11082, 72.98961, 73.16777, 73.36272, 73.0228, 71.28471,
  93.37275, 93.91972, 94.21539, 94.34156, 94.75257, 95.10362, 95.4132, 
    95.79151, 94.46622, 94.86961, 95.07227, 95.66429, 95.79955, 95.95409, 
    96.39525, 96.7307, 95.6562, 95.84826, 96.22713, 96.19344,
  88.12901, 88.89231, 89.7457, 90.62141, 91.49396, 92.44537, 93.39051, 
    94.25302, 91.01757, 91.81031, 92.62436, 93.2332, 93.95383, 94.29411, 
    94.67218, 94.90065, 93.31431, 94.06856, 94.98056, 95.90086,
  87.34212, 89.01546, 90.59021, 92.04594, 93.36865, 94.53568, 95.52061, 
    96.28748, 91.86085, 92.71123, 93.42807, 94.01946, 94.74444, 95.34738, 
    95.41664, 96.01217, 94.65759, 95.64129, 96.25311, 96.99723,
  86.33559, 88.1441, 89.5666, 91.11248, 92.25186, 93.53372, 94.53056, 
    95.21667, 92.55618, 93.30819, 94.12542, 94.77509, 95.55293, 96.51119, 
    97.34533, 97.95737, 98.86752, 99.07931, 98.6409, 98.26416,
  84.34882, 85.62908, 86.99768, 87.90079, 88.35789, 88.64817, 89.12117, 
    90.08427, 89.70327, 90.78755, 91.51633, 90.93925, 91.52043, 92.58109, 
    93.84431, 94.75764, 97.23259, 97.36762, 97.09634, 96.73912,
  83.37933, 85.54396, 86.65485, 87.35948, 88.15724, 88.7373, 89.02234, 
    89.13257, 84.65704, 85.29153, 85.96129, 86.39213, 86.97983, 87.81332, 
    88.90668, 89.84061, 95.99057, 96.46244, 95.87488, 95.04823,
  91.26807, 90.90514, 91.1543, 90.93425, 91.22235, 92.76355, 92.37339, 
    91.95372, 84.30848, 83.99349, 84.40256, 80.3712, 81.53752, 86.64213, 
    90.45585, 87.53249, 92.90964, 94.03133, 94.93694, 95.31119,
  71.14718, 69.40942, 67.96175, 66.10277, 67.23072, 69.91323, 68.59761, 
    66.8392, 61.88372, 64.66482, 72.10359, 79.0449, 81.94794, 87.70512, 
    91.49586, 91.20327, 93.17608, 92.24327, 90.30618, 89.61055,
  69.44691, 67.61513, 66.10161, 65.21225, 64.9798, 65.75106, 67.18806, 
    68.39124, 67.0039, 67.0452, 66.92162, 68.55112, 72.37344, 76.01417, 
    79.56667, 82.39173, 85.5618, 89.72083, 90.78975, 93.5921,
  76.7655, 76.04768, 75.18473, 74.02251, 73.11304, 73.20016, 74.07021, 
    74.83585, 75.77511, 76.08671, 76.19196, 76.03816, 75.69469, 75.63595, 
    75.73514, 76.87009, 79.41619, 82.42207, 84.44841, 85.53425,
  82.92245, 82.35838, 81.8168, 80.87459, 79.7678, 79.37811, 79.88898, 
    81.15392, 82.12207, 81.77625, 81.58807, 81.76734, 81.67142, 81.26604, 
    81.16002, 81.75224, 82.56812, 82.80696, 82.80157, 83.63928,
  85.94359, 86.2039, 86.42712, 86.53812, 85.87373, 84.22209, 82.8445, 
    83.56202, 85.77419, 86.76926, 86.77412, 86.74758, 86.60226, 86.6552, 
    86.95509, 86.90311, 86.93803, 86.04026, 83.97957, 82.545,
  86.72565, 87.57019, 87.79339, 88.12904, 87.90759, 85.7135, 82.6209, 
    80.8781, 81.59084, 83.24759, 85.08566, 86.95364, 88.3853, 88.82724, 
    89.19962, 89.26579, 88.1617, 86.47892, 84.71124, 82.30123,
  82.75827, 82.88097, 82.8921, 82.43293, 81.3303, 79.89459, 78.65818, 78.202, 
    78.84344, 80.26993, 82.08205, 84.45817, 86.92677, 88.15726, 88.65891, 
    88.66456, 86.91369, 85.5312, 85.49545, 84.94057,
  78.13414, 76.37182, 76.15897, 76.39225, 75.88791, 75.69257, 76.51527, 
    78.30303, 80.59325, 83.04788, 85.2299, 87.10377, 88.48997, 88.60088, 
    88.72065, 89.11111, 88.57193, 87.63721, 87.81053, 88.19389,
  73.66436, 72.32921, 72.67623, 74.37872, 75.73877, 77.11079, 78.95532, 
    81.16214, 83.66551, 85.66153, 87.16323, 88.23895, 89.21335, 89.94067, 
    90.56502, 90.74302, 90.11922, 89.17405, 89.16929, 88.38626,
  71.18357, 72.14453, 74.02247, 75.90031, 77.01978, 78.2691, 79.49795, 
    79.92043, 80.67075, 82.46883, 84.50685, 86.37706, 87.82352, 88.65002, 
    89.12348, 89.50642, 88.54946, 86.60401, 85.23292, 83.90275,
  73.10514, 74.22552, 75.39771, 76.09384, 76.31498, 76.84937, 76.481, 
    73.56741, 70.80209, 72.01581, 75.74261, 79.66776, 82.23591, 83.46809, 
    84.10751, 84.67477, 82.85084, 79.45297, 77.64763, 77.45921,
  74.51862, 74.8261, 73.29723, 71.60673, 71.36654, 72.10418, 70.09155, 
    66.58561, 64.47836, 64.06046, 65.22453, 68.07657, 71.73197, 74.37994, 
    75.76649, 75.4369, 73.96723, 73.12037, 74.10836, 75.17548,
  71.20527, 69.69956, 66.79221, 65.56136, 68.20262, 69.70413, 69.78534, 
    68.38866, 69.32178, 69.11639, 66.99824, 67.11583, 70.60143, 74.46976, 
    75.0638, 73.81257, 73.84793, 75.27972, 76.86605, 76.99019,
  90.07456, 90.48672, 90.86421, 91.27199, 91.64136, 92.08289, 92.41364, 
    92.75996, 91.4425, 91.91649, 92.32284, 92.60006, 92.81592, 93.39871, 
    93.97868, 94.02592, 93.36269, 93.66527, 94.14593, 94.19774,
  84.29382, 85.41369, 86.9097, 88.23539, 89.8544, 91.51548, 92.97314, 
    94.33192, 91.55229, 92.75607, 93.37475, 94.15374, 94.3779, 94.60982, 
    94.75601, 95.42723, 93.769, 95.04896, 95.64101, 97.12575,
  86.82552, 88.53922, 90.2179, 91.6937, 92.82541, 93.79211, 94.62707, 
    95.27658, 90.75754, 92.08592, 93.7529, 95.66997, 96.54538, 96.90233, 
    96.83202, 96.85136, 96.48665, 97.25517, 97.1412, 97.36676,
  86.51781, 88.45362, 90.30604, 91.7568, 93.23621, 94.36797, 94.71826, 
    94.96798, 93.05251, 94.24355, 95.3751, 96.8235, 98.503, 99.18272, 
    99.18351, 99.02308, 98.74769, 98.01578, 97.30558, 96.38832,
  84.19908, 86.45179, 88.48095, 89.98982, 90.51294, 90.4688, 90.82926, 
    91.86302, 91.82877, 93.24203, 94.43957, 94.97415, 95.24644, 96.79502, 
    98.19026, 98.66412, 99.60326, 99.62563, 99.20312, 98.10313,
  84.45502, 84.94581, 86.16518, 87.34177, 87.47768, 86.88894, 86.37795, 
    86.30563, 82.23832, 82.71339, 83.38699, 83.94523, 85.16924, 86.55328, 
    87.96186, 89.21535, 95.08026, 95.72395, 96.02077, 96.26938,
  95.16702, 92.33752, 90.27086, 89.07218, 88.38104, 88.88416, 89.29356, 
    90.25732, 83.33585, 84.71282, 86.10643, 80.853, 83.1026, 88.52948, 
    91.32358, 87.85949, 92.61178, 93.57198, 94.85641, 95.65263,
  90.04991, 87.42262, 84.45006, 83.09418, 82.52718, 84.89194, 87.55519, 
    89.00037, 83.30129, 85.12016, 88.76704, 87.65919, 88.64612, 91.80663, 
    95.6026, 96.06413, 96.26199, 95.8017, 95.25934, 95.15553,
  71.42123, 69.97279, 68.28963, 66.32768, 65.43402, 65.7264, 66.14357, 
    67.20413, 67.14657, 68.20274, 71.70902, 76.28211, 81.89819, 85.73148, 
    87.89687, 89.7194, 92.84814, 94.96597, 96.06687, 95.8121,
  78.0134, 78.29984, 77.96667, 76.92651, 75.44479, 74.00323, 73.11319, 
    72.67534, 72.69421, 72.11981, 71.96851, 72.5605, 72.955, 72.42447, 
    71.92396, 71.87505, 71.97475, 73.14788, 75.44102, 77.93836,
  85.37109, 85.71864, 85.34331, 84.56796, 83.66139, 82.60973, 81.97827, 
    81.90745, 82.00715, 81.58857, 81.45783, 81.49622, 81.26762, 80.44291, 
    79.70499, 78.92028, 77.4854, 75.70467, 74.76763, 75.75611,
  87.15807, 87.70086, 87.97696, 88.21327, 88.03773, 86.19876, 84.38065, 
    84.94342, 87.52986, 88.90504, 88.68471, 87.89834, 86.94041, 86.22071, 
    85.76936, 84.88177, 83.09745, 80.65755, 77.76865, 76.11965,
  85.23028, 86.15197, 86.90668, 88.18147, 89.40193, 88.46203, 85.715, 
    83.90537, 84.75997, 86.61617, 87.65101, 88.08749, 88.34624, 88.50468, 
    88.86424, 88.98323, 87.28278, 84.29656, 81.63602, 79.26149,
  82.01743, 82.46607, 83.36809, 84.53693, 84.61572, 83.5394, 82.01644, 
    81.28974, 82.30324, 83.89819, 85.27593, 86.587, 87.77227, 88.66557, 
    89.16769, 89.02431, 87.08436, 85.04607, 84.15939, 83.59784,
  78.719, 76.68517, 76.54944, 77.59534, 77.64058, 77.25024, 77.12875, 
    78.08372, 80.3743, 82.90988, 85.57194, 87.5092, 88.51685, 88.79141, 
    88.48484, 87.72935, 86.21063, 84.72538, 85.0446, 85.67335,
  72.91538, 70.91225, 70.40004, 72.00016, 73.97049, 75.86927, 78.27828, 
    81.14394, 83.91167, 86.30752, 88.2465, 89.2392, 89.80845, 89.84117, 
    88.67654, 87.81126, 86.84928, 85.75919, 85.76432, 84.81652,
  68.98612, 70.11836, 72.07506, 74.48186, 76.79041, 78.84361, 80.78701, 
    82.70566, 84.8105, 87.28165, 88.81762, 89.28561, 89.12044, 88.63956, 
    87.3147, 86.41982, 85.03951, 83.22682, 81.85175, 80.65599,
  71.87428, 73.88077, 75.56699, 76.5269, 77.06773, 78.18127, 78.06432, 
    74.25318, 71.11487, 72.67726, 76.20137, 79.51053, 81.47756, 81.98953, 
    81.87717, 81.5437, 79.3908, 76.54128, 74.65981, 74.18701,
  71.2946, 71.91714, 71.57894, 70.90557, 71.9691, 72.63856, 68.89857, 
    64.0445, 62.01991, 61.49824, 62.49363, 64.22562, 67.11063, 69.33882, 
    70.72939, 71.53349, 71.32391, 70.3533, 70.42554, 72.01726,
  65.94721, 65.21111, 64.98637, 66.46193, 69.14471, 69.29983, 69.35908, 
    67.34663, 69.33524, 69.58876, 65.63332, 64.47161, 68.88573, 72.17902, 
    72.74658, 73.30175, 73.66959, 73.32896, 72.45762, 71.98344,
  91.17011, 91.58001, 91.85252, 92.27715, 92.66914, 93.01484, 93.47704, 
    93.82074, 92.58183, 93.19258, 93.38977, 93.6412, 94.05588, 94.41631, 
    94.68109, 94.93601, 94.35142, 94.49462, 94.546, 94.59042,
  86.77498, 88.07269, 89.27798, 90.34485, 91.55575, 92.46603, 93.63637, 
    94.69076, 91.81561, 92.89853, 93.56634, 94.50151, 95.24194, 96.23975, 
    97.06346, 97.78746, 96.53555, 96.97373, 97.45118, 97.49062,
  86.59285, 88.4179, 90.03355, 91.04927, 91.9567, 92.99967, 94.0715, 
    94.96685, 91.05003, 92.6053, 94.1451, 95.61274, 96.81329, 97.89839, 
    98.22961, 98.41768, 98.01109, 98.2739, 98.72503, 99.02295,
  85.72983, 87.67071, 89.67376, 91.36398, 92.63693, 93.82869, 94.73441, 
    96.05701, 94.43509, 95.67455, 96.84856, 97.83617, 98.55512, 99.01227, 
    99.24763, 99.30426, 98.92216, 98.3271, 98.91103, 99.14411,
  83.84087, 85.55367, 86.6799, 88.35298, 90.05916, 91.30825, 92.77764, 
    94.5013, 95.06129, 96.50959, 97.56435, 98.22564, 98.49876, 98.56296, 
    98.71836, 98.61203, 99.80033, 99.65018, 99.5316, 99.62746,
  81.29015, 82.9984, 84.57397, 86.78717, 88.33836, 89.20285, 89.8382, 
    90.01332, 86.25098, 86.94479, 87.62567, 88.50341, 89.89535, 91.3922, 
    92.65845, 93.59153, 98.44129, 98.56503, 98.68295, 98.1797,
  94.11578, 89.39543, 88.14638, 88.23101, 88.19188, 88.5246, 88.8085, 
    89.19108, 81.55666, 81.38972, 82.86344, 78.6693, 80.35023, 86.70567, 
    89.25298, 89.13045, 94.88373, 95.91883, 96.15907, 95.86631,
  93.47617, 93.4659, 93.94927, 94.54108, 94.8801, 96.0095, 96.58344, 
    96.88368, 94.05307, 93.64865, 95.48979, 92.48824, 92.40602, 94.77396, 
    96.82478, 97.08608, 97.73698, 97.53609, 93.8558, 93.96168,
  85.90707, 86.48092, 88.41611, 90.64163, 91.81621, 92.8755, 94.00491, 
    95.20415, 94.20609, 94.29536, 94.39256, 94.48383, 95.0556, 95.36298, 
    95.81496, 95.94225, 97.36671, 98.47647, 98.54305, 96.72159,
  72.88133, 74.20032, 74.76454, 76.1488, 77.4093, 79.06323, 81.18011, 
    83.68102, 85.68005, 85.24361, 84.31608, 84.50407, 85.39473, 84.996, 
    84.42863, 85.12097, 86.13593, 88.14323, 90.67519, 93.00241,
  66.63493, 68.23456, 67.53545, 65.99398, 65.89098, 65.93284, 66.67316, 
    68.94611, 71.95542, 72.95057, 73.88634, 75.06085, 76.0082, 76.36845, 
    76.31053, 75.89989, 75.37329, 74.22463, 73.36652, 73.20379,
  69.53298, 71.56736, 73.28878, 74.78682, 75.60504, 74.75257, 73.83785, 
    74.73756, 78.06574, 80.53299, 81.91823, 82.66595, 82.96272, 83.04848, 
    82.81315, 82.33181, 81.64347, 80.23748, 78.04977, 76.26704,
  74.75862, 76.4924, 77.82009, 79.74557, 81.41613, 81.71525, 80.41744, 
    79.33185, 80.11401, 81.40411, 82.73872, 83.85191, 84.49371, 84.17726, 
    84.05972, 84.38174, 83.88985, 82.7181, 81.48486, 80.10326,
  73.93359, 74.53183, 75.94057, 77.88861, 79.19852, 79.60794, 79.20315, 
    78.43513, 78.54962, 79.61915, 81.24841, 82.89156, 84.24147, 85.2039, 
    86.23164, 86.99693, 85.79055, 84.85445, 84.519, 84.11481,
  71.76712, 70.07494, 70.63139, 72.36175, 73.28513, 74.11209, 75.00201, 
    75.93827, 78.47118, 81.37273, 84.69566, 87.34113, 88.61317, 89.30084, 
    89.70651, 89.7278, 88.04289, 86.20798, 85.52447, 85.30213,
  66.02827, 64.54211, 64.65984, 66.86544, 69.47443, 72.26003, 75.21101, 
    78.47057, 82.4762, 85.68998, 88.68793, 90.65517, 91.84777, 92.5185, 
    92.34897, 91.22189, 89.04608, 86.93361, 86.25781, 85.16582,
  61.84498, 63.78832, 66.99315, 70.68969, 73.75171, 76.79504, 79.40872, 
    81.17258, 83.29347, 85.87012, 88.92642, 91.04924, 91.7319, 92.00223, 
    91.74808, 90.20827, 88.03146, 85.93414, 84.358, 83.12246,
  67.2907, 70.96338, 74.56693, 76.99506, 77.73013, 78.31666, 77.02131, 
    71.61569, 69.24093, 71.21501, 76.57626, 82.15186, 85.38359, 86.74759, 
    86.68133, 85.62526, 82.71592, 78.63671, 75.73563, 74.57832,
  73.94997, 76.4595, 77.19582, 75.5669, 74.13396, 71.82111, 65.86146, 
    61.56705, 61.72529, 61.04848, 62.0101, 65.11713, 70.12402, 72.49516, 
    71.98722, 70.99656, 69.32114, 67.64272, 67.41056, 68.16187,
  73.51095, 72.88679, 70.64802, 68.74767, 69.36805, 67.2804, 65.18354, 
    62.87301, 64.75318, 65.11667, 61.41754, 62.05071, 68.23034, 72.16243, 
    71.34657, 70.70106, 69.99625, 69.40432, 69.33576, 68.67924,
  90.98745, 91.29696, 91.60209, 92.00352, 92.26562, 92.61909, 93.00459, 
    93.36853, 92.07767, 92.36163, 92.46584, 92.6298, 93.01018, 93.3162, 
    93.62531, 94.05055, 93.27223, 93.43857, 93.69898, 93.74854,
  85.01886, 86.37234, 87.72834, 89.1521, 90.49723, 91.81866, 92.91039, 
    94.00024, 90.70879, 91.43392, 91.81021, 91.96034, 92.56762, 93.55199, 
    94.66047, 95.84389, 94.8726, 95.92691, 96.81916, 97.21001,
  83.95771, 86.06379, 88.0361, 89.80649, 91.38123, 92.52282, 93.28365, 
    93.86976, 89.2356, 90.37859, 92.15395, 93.23993, 94.22323, 95.09611, 
    96.2742, 97.27421, 96.27925, 96.46619, 96.57714, 96.53323,
  85.6008, 87.56618, 89.47357, 91.66181, 93.33055, 94.50098, 95.13374, 
    94.89646, 92.98121, 94.14777, 95.11217, 96.46093, 97.58001, 98.52686, 
    99.29742, 99.38843, 99.58778, 99.05384, 98.16373, 97.20988,
  85.5621, 88.19527, 90.44502, 91.62866, 91.73222, 92.1685, 92.03563, 
    92.00865, 91.9073, 92.9025, 93.7832, 94.50246, 95.14792, 95.83698, 
    96.59937, 97.10381, 99.25783, 99.54443, 99.38344, 98.83322,
  84.65897, 86.63267, 87.36778, 88.36446, 88.97176, 89.78, 90.15521, 
    90.34492, 86.21194, 86.44642, 87.18334, 88.40533, 89.90788, 91.47908, 
    92.76173, 93.2648, 97.67901, 97.69427, 97.95529, 98.23748,
  93.90025, 92.46072, 92.43479, 92.6404, 92.80974, 93.12684, 93.19376, 
    92.79742, 84.05801, 84.57143, 86.53767, 83.70232, 85.1542, 88.3131, 
    89.87689, 88.88409, 92.52689, 92.21806, 92.1344, 91.90836,
  96.93919, 97.68593, 97.96864, 97.89955, 97.66016, 97.79575, 97.30118, 
    96.62569, 91.55299, 91.37716, 92.15118, 87.67492, 88.36038, 90.62241, 
    93.78268, 94.54948, 95.53249, 95.10094, 91.58355, 91.0564,
  98.32555, 97.83466, 97.6034, 97.96844, 98.39095, 98.83584, 98.88914, 
    98.20824, 96.4235, 96.60486, 96.46543, 96.09408, 95.59052, 94.93619, 
    94.23808, 94.4162, 95.42523, 96.56586, 96.63497, 95.78254,
  98.12569, 98.27222, 97.82526, 97.16116, 96.27717, 95.64143, 95.25061, 
    95.17387, 95.88683, 96.99593, 98.4914, 99.04877, 99.34573, 99.13908, 
    98.3607, 96.95287, 95.44658, 93.61249, 93.62886, 95.46103,
  94.96774, 95.5589, 95.26688, 93.56842, 87.32948, 82.36816, 83.5425, 
    89.27451, 92.10559, 92.78727, 92.4663, 91.67569, 89.4976, 87.5445, 
    86.24968, 82.81287, 76.93233, 74.39601, 74.04531, 75.7169,
  72.37726, 73.68614, 72.95264, 70.60884, 64.085, 58.66286, 57.24234, 
    59.58153, 64.93045, 68.80866, 70.19659, 70.7561, 72.11375, 74.55909, 
    77.05973, 77.96165, 78.4235, 77.22953, 74.56795, 73.03501,
  60.79295, 62.42181, 63.15622, 63.12088, 62.95715, 62.28113, 61.18781, 
    61.19473, 62.61267, 64.99561, 67.12331, 69.33784, 72.38282, 76.10181, 
    80.3075, 82.50353, 83.20199, 81.96946, 80.01646, 78.29514,
  62.52289, 62.34185, 62.01292, 61.60038, 61.29708, 61.24829, 61.4658, 
    61.92487, 62.66392, 63.96798, 65.79452, 69.01866, 73.35307, 78.09818, 
    82.1577, 84.98119, 85.99424, 85.79336, 85.78348, 85.27866,
  63.34808, 60.43627, 58.75488, 58.37927, 58.04855, 58.33051, 59.3683, 
    60.48534, 62.1982, 64.82623, 68.62986, 73.79235, 78.38273, 81.82935, 
    84.18407, 85.44627, 85.53128, 84.86642, 85.29137, 86.35084,
  62.13792, 58.48501, 56.34128, 56.65401, 58.03448, 59.82373, 61.8807, 
    64.58637, 68.92142, 73.62315, 77.8894, 81.73029, 84.82333, 86.50983, 
    86.46868, 85.33784, 84.00378, 83.01505, 83.86026, 84.7075,
  58.99577, 58.11288, 59.93508, 63.42055, 66.57792, 69.12582, 71.43848, 
    73.48515, 76.22089, 79.1198, 81.74926, 83.83871, 85.40308, 86.47977, 
    86.28207, 85.2745, 83.37839, 81.258, 80.58562, 80.90097,
  63.8393, 67.91364, 72.20181, 74.81266, 75.83478, 76.13286, 73.61414, 
    68.05742, 65.72118, 66.67308, 69.43307, 72.90327, 76.30459, 78.75282, 
    80.40519, 80.60797, 77.91299, 73.88861, 71.77665, 71.94137,
  71.71375, 74.3072, 75.18604, 74.75976, 75.20363, 72.63457, 65.05898, 
    60.53121, 59.03997, 56.64069, 55.9188, 57.47602, 60.75026, 64.24229, 
    66.50427, 67.12095, 66.49196, 66.05244, 67.14204, 69.58089,
  69.12215, 69.33967, 68.79024, 69.13474, 71.21356, 68.23521, 65.90282, 
    65.22256, 64.527, 61.75634, 57.16112, 57.24561, 62.23014, 66.12975, 
    67.02992, 67.16248, 68.56287, 71.1139, 74.02827, 75.82978,
  92.8159, 93.2197, 93.6105, 93.91306, 94.22326, 94.58191, 94.92522, 
    95.22913, 93.85856, 94.2981, 94.47391, 94.7088, 95.17386, 95.4691, 
    95.4802, 95.73299, 95.02055, 95.20663, 95.11687, 95.06095,
  86.55241, 87.79284, 89.09595, 90.32372, 91.73504, 93.10539, 94.27875, 
    95.06039, 91.63329, 92.67184, 93.37179, 93.94209, 94.32087, 95.02787, 
    95.71693, 96.00041, 94.48289, 95.29887, 96.84354, 97.49466,
  85.51675, 86.73094, 88.12775, 89.64433, 91.18484, 92.60871, 94.02316, 
    95.21175, 90.87081, 92.2225, 92.91127, 94.14934, 94.48235, 95.27862, 
    95.96638, 96.41363, 96.01525, 96.78755, 97.30156, 97.7453,
  87.86299, 89.97968, 91.36497, 92.4736, 93.3867, 94.78036, 96.14001, 
    97.43903, 95.68842, 97.21931, 98.24479, 98.87528, 99.1653, 99.05997, 
    99.26906, 99.32961, 99.47722, 99.5089, 99.29516, 99.02122,
  83.55333, 86.24703, 88.14996, 90.44866, 92.48737, 94.4408, 95.76079, 
    96.25528, 95.86619, 96.43434, 96.67438, 96.65849, 96.37702, 96.32846, 
    96.70243, 96.93121, 98.8772, 98.80267, 98.70007, 98.47133,
  82.02061, 83.96915, 85.86088, 87.45531, 88.73535, 89.68233, 89.84081, 
    89.59205, 85.68663, 86.62338, 87.67474, 88.7756, 89.80199, 90.61549, 
    91.45695, 92.18902, 97.42504, 97.88176, 98.10278, 97.82326,
  94.65263, 91.70213, 91.08222, 90.87824, 90.92789, 91.0863, 89.85123, 
    88.96008, 79.85953, 79.76646, 81.62791, 78.33206, 80.6271, 86.04789, 
    88.08054, 88.24763, 93.84735, 94.6907, 95.16203, 94.95577,
  98.42578, 98.40656, 98.55572, 97.96102, 97.41238, 97.13661, 96.55749, 
    96.29939, 91.6566, 91.80348, 92.40903, 89.13735, 89.5166, 92.98286, 
    95.18192, 92.46988, 95.14555, 94.10226, 93.30116, 93.54501,
  97.54238, 97.18066, 96.43796, 95.75636, 95.22883, 95.55516, 96.3735, 
    97.04151, 95.48612, 95.69362, 95.47098, 95.28168, 94.99551, 94.68185, 
    95.20041, 96.02824, 96.93748, 97.56205, 97.4871, 97.27131,
  95.49395, 95.33186, 94.76794, 93.87866, 93.72905, 93.85388, 93.78401, 
    94.40219, 95.28983, 96.78725, 97.46341, 98.35218, 98.66293, 98.68405, 
    98.70512, 98.38976, 97.50048, 96.24825, 96.30229, 96.65794,
  96.56091, 96.8774, 96.98513, 96.51257, 95.94294, 94.89609, 94.397, 
    94.50034, 95.31358, 95.6545, 96.15311, 96.7962, 96.82693, 96.65706, 
    96.53819, 94.64299, 87.44152, 72.86719, 67.6725, 70.70515,
  93.95828, 93.95774, 93.69702, 93.56377, 92.41996, 81.67066, 72.72379, 
    69.24843, 73.34854, 80.0995, 82.82, 81.80415, 79.01461, 76.48002, 
    75.28624, 72.49391, 69.0419, 65.5322, 63.06635, 62.98507,
  75.39345, 75.21915, 74.39631, 74.04247, 73.37346, 69.44512, 64.82233, 
    62.41673, 62.08951, 62.96581, 63.79028, 64.37586, 64.81615, 65.71603, 
    68.6466, 70.66341, 71.33911, 70.47929, 68.89828, 68.01688,
  72.86983, 71.53578, 70.28037, 69.1014, 67.61387, 66.09517, 64.6434, 
    63.52663, 63.60285, 64.69032, 65.69706, 67.03696, 69.1563, 71.72166, 
    73.77777, 75.05098, 74.70728, 74.41285, 74.35855, 74.02293,
  73.2523, 69.52663, 66.16081, 63.94156, 61.83159, 60.53927, 60.05917, 
    60.40867, 61.74479, 63.5501, 65.86928, 68.87156, 72.5392, 75.67437, 
    77.1875, 77.49569, 76.67693, 75.47895, 75.01425, 75.11897,
  70.58049, 66.28109, 62.42197, 61.03706, 60.57674, 60.737, 61.45941, 
    62.96795, 65.5925, 69.01488, 72.80242, 76.15392, 78.67603, 80.11696, 
    80.21175, 79.41575, 77.46162, 75.06468, 74.20818, 73.83661,
  63.8953, 62.55087, 63.60147, 66.0998, 67.4076, 68.06668, 68.99622, 
    70.18645, 71.72113, 74.77647, 78.03604, 80.17949, 81.32273, 81.70218, 
    81.14687, 79.72179, 76.58879, 73.3121, 71.03906, 70.11959,
  65.15434, 69.2553, 74.13488, 76.44986, 76.32185, 74.95175, 71.48375, 
    65.98779, 62.8257, 63.31886, 66.21056, 69.7999, 72.91084, 75.24597, 
    76.60191, 75.72329, 71.19488, 65.76025, 62.80171, 61.90194,
  76.43947, 79.50707, 80.23241, 77.65983, 74.37008, 69.15773, 61.65321, 
    57.76416, 56.00876, 53.5259, 52.2877, 53.15834, 55.19382, 58.31443, 
    61.5801, 62.28934, 61.09306, 59.53255, 59.20259, 59.69647,
  78.29018, 77.09428, 74.13283, 70.94929, 69.28881, 64.00248, 61.85705, 
    64.93412, 63.97273, 60.72979, 54.75216, 54.21546, 58.42363, 62.03396, 
    63.6741, 64.19766, 64.62788, 65.13469, 65.96899, 66.69779,
  93.69763, 93.98157, 94.17415, 94.62468, 94.92327, 95.37312, 95.63943, 
    95.98896, 94.81039, 95.14245, 95.41955, 95.74541, 96.00251, 96.22443, 
    96.50529, 96.65051, 96.10497, 96.03961, 96.41432, 96.76353,
  88.61023, 89.30877, 89.85851, 90.45193, 91.32699, 92.22941, 93.21968, 
    94.25391, 91.21249, 92.17634, 93.1927, 94.04564, 94.70544, 95.26926, 
    95.60767, 96.08686, 94.31548, 94.89679, 95.44227, 95.96345,
  85.20106, 86.95082, 88.75328, 90.41666, 92.0328, 93.31853, 94.25261, 
    95.16662, 91.08914, 92.01147, 92.61927, 93.14661, 94.26891, 95.15186, 
    95.31612, 95.59884, 94.56198, 95.1679, 95.89069, 96.52539,
  87.37148, 89.41404, 90.92465, 91.76102, 92.70269, 93.31511, 93.52556, 
    94.36659, 92.01796, 93.38969, 94.90091, 95.91694, 96.57777, 97.30638, 
    97.93712, 98.58411, 99.34196, 99.7229, 99.80676, 99.27079,
  84.38491, 86.47743, 88.5022, 89.71974, 90.95544, 92.29185, 93.52992, 
    94.20676, 93.95078, 94.43997, 94.26513, 93.72448, 93.66109, 94.52975, 
    95.29276, 96.14672, 98.62106, 99.02883, 99.11876, 99.1041,
  82.98889, 84.79034, 85.99445, 87.29128, 88.4016, 89.1859, 90.24387, 
    90.87609, 86.84308, 86.65687, 86.22065, 86.9841, 88.03822, 89.34309, 
    90.55196, 91.74538, 97.54018, 98.22718, 98.55006, 97.86477,
  95.70589, 92.68562, 92.32629, 92.23976, 91.71163, 91.91738, 91.75796, 
    91.22165, 82.03094, 81.57092, 82.16418, 77.62531, 78.72924, 84.20027, 
    85.59505, 83.81256, 90.85746, 92.08733, 93.0552, 93.16888,
  99.13496, 99.54393, 99.4279, 98.80517, 98.187, 98.37833, 98.96397, 
    99.22973, 95.61932, 95.84886, 96.04897, 94.25564, 94.14145, 95.16939, 
    94.79033, 90.53915, 93.59682, 92.63699, 88.32133, 88.61066,
  98.32017, 98.91051, 99.14117, 99.07484, 99.04048, 98.96371, 98.63768, 
    98.62859, 97.90269, 98.24556, 98.49007, 98.75141, 98.4716, 97.96627, 
    97.89454, 97.48149, 97.28754, 97.66056, 97.0302, 96.41569,
  96.73216, 97.23348, 97.65511, 97.85133, 98.05978, 97.95016, 97.74843, 
    97.82138, 97.88368, 97.39843, 96.52958, 96.88121, 96.51434, 96.92643, 
    98.12704, 98.42097, 97.91376, 97.33286, 97.05994, 96.59552,
  96.0761, 96.68906, 97.18467, 97.16145, 97.49075, 96.83777, 96.40249, 
    97.06275, 97.23053, 96.84941, 96.53326, 96.5626, 96.82115, 95.80025, 
    95.65185, 96.09574, 95.88062, 92.6073, 85.5697, 80.2245,
  96.28162, 95.91197, 95.11305, 95.37505, 96.24417, 93.95023, 86.0817, 
    79.15984, 78.62903, 84.00212, 90.78424, 92.53625, 91.86491, 90.9398, 
    92.07838, 91.50728, 87.51357, 77.07855, 65.62537, 58.9409,
  77.90456, 77.93506, 78.87369, 78.57576, 78.47137, 74.99793, 67.78358, 
    62.05617, 61.52721, 63.17921, 64.6997, 65.4013, 65.71869, 66.27252, 
    67.61083, 69.40225, 69.7475, 67.13508, 63.55815, 62.26278,
  69.71602, 68.81417, 67.97478, 67.09431, 65.83036, 64.0762, 62.32809, 
    61.61483, 61.742, 63.08266, 64.50009, 66.0673, 67.9017, 70.04298, 
    72.29219, 74.09147, 73.16489, 72.29854, 71.26584, 69.51695,
  69.65104, 66.6459, 64.56651, 63.05555, 61.35976, 59.80534, 59.00587, 
    59.22359, 60.82201, 63.74959, 66.91178, 69.95277, 72.88194, 75.39922, 
    77.28359, 78.3858, 77.79736, 76.7859, 75.90878, 75.02176,
  66.45039, 62.7214, 58.99157, 57.04194, 56.59826, 57.54989, 59.27354, 
    62.10122, 66.43124, 70.93253, 74.74186, 77.98203, 80.50579, 82.1219, 
    82.28754, 81.49641, 79.55513, 77.50551, 76.76811, 75.89095,
  59.8067, 57.19482, 56.45367, 57.96009, 59.69281, 61.96859, 65.10448, 
    68.9625, 73.21517, 76.74874, 79.04732, 80.4557, 81.70774, 82.91959, 
    82.80328, 81.73381, 79.18402, 76.22301, 73.41568, 71.17374,
  62.50906, 64.62785, 67.70721, 70.20687, 71.38424, 72.12524, 71.30563, 
    68.77511, 66.99574, 67.47031, 69.20536, 71.10355, 73.62134, 75.74953, 
    76.93594, 76.81344, 73.34011, 68.27863, 64.62132, 62.55026,
  74.45332, 77.16498, 77.91454, 77.22263, 76.25582, 72.94933, 67.16231, 
    64.12454, 62.84193, 60.16876, 58.80754, 59.71167, 61.71157, 63.64535, 
    65.34641, 65.56149, 64.05979, 62.48677, 62.16053, 62.83937,
  76.36472, 76.32736, 75.03173, 73.49324, 72.97213, 68.37362, 66.42924, 
    68.67296, 69.40749, 67.33298, 62.51077, 62.30519, 67.18233, 68.27329, 
    67.70455, 67.42226, 67.46717, 67.80292, 69.4464, 71.91476,
  93.0022, 93.54292, 93.79911, 94.09368, 94.70123, 95.14903, 95.5219, 
    95.85071, 94.32282, 94.82507, 95.2749, 95.55389, 95.9054, 96.1316, 
    96.46326, 96.78541, 96.08192, 96.39866, 96.39725, 96.78385,
  85.02152, 86.42142, 87.75742, 89.28708, 90.6942, 92.29068, 93.56042, 
    94.86628, 91.66965, 92.96471, 93.56914, 94.88222, 95.54645, 96.09328, 
    96.35301, 96.64264, 95.26493, 96.02611, 96.3009, 97.1591,
  82.62967, 85.39384, 88.17564, 90.64791, 92.49731, 93.85115, 94.84271, 
    95.74956, 91.06268, 92.37741, 93.46746, 95.01662, 96.24152, 97.20704, 
    98.19744, 99.11477, 98.84184, 99.33872, 99.42726, 99.59704,
  85.38585, 87.92935, 90.29302, 92.16904, 93.91631, 95.36686, 96.41099, 
    97.22126, 95.25395, 96.47607, 97.69157, 98.55507, 99.24526, 99.58598, 
    99.72582, 99.76407, 99.89597, 99.86573, 99.83057, 99.67528,
  82.96909, 85.34504, 87.31969, 89.28407, 91.31425, 93.1142, 93.89056, 
    94.04408, 93.53922, 93.97161, 94.85207, 95.86453, 96.87653, 97.549, 
    98.06141, 98.71509, 99.9036, 99.96779, 99.72726, 99.1424,
  79.42523, 81.14129, 82.46816, 83.58894, 84.28524, 84.70596, 85.89222, 
    87.56048, 84.54214, 85.79517, 87.01311, 88.1989, 89.20309, 90.33458, 
    91.0071, 91.93439, 96.75284, 97.07966, 97.19107, 96.92353,
  93.06845, 91.78378, 90.74979, 89.19584, 88.54763, 88.41358, 88.77499, 
    89.38712, 81.95401, 82.87835, 85.87792, 77.2277, 78.48421, 85.97547, 
    87.55101, 83.68902, 89.86437, 91.42082, 92.65909, 93.37128,
  96.98489, 97.29073, 96.91201, 95.66315, 95.45506, 95.88181, 96.86057, 
    97.46348, 94.02431, 94.93224, 96.48778, 92.778, 93.11106, 96.12519, 
    98.01921, 90.32995, 96.12097, 93.41193, 89.77426, 90.8561,
  97.73721, 97.65613, 97.70346, 97.68906, 97.49747, 97.26411, 97.00942, 
    96.75341, 95.36272, 95.82192, 96.45075, 96.55427, 96.61069, 96.8299, 
    97.13477, 97.74607, 98.52603, 99.11051, 98.78793, 98.49687,
  95.51378, 95.65935, 95.6003, 95.42876, 95.931, 96.26857, 96.15498, 96.2915, 
    96.63461, 96.92522, 96.99387, 96.94753, 97.21856, 96.79762, 96.9921, 
    97.44846, 97.49514, 97.34497, 97.28771, 96.9775,
  95.03127, 95.21569, 95.30614, 95.11676, 94.97446, 94.78693, 94.78231, 
    94.94573, 95.57629, 96.11303, 96.05106, 95.87893, 95.45326, 95.0597, 
    95.02916, 94.73145, 93.87691, 93.1442, 91.39059, 89.31501,
  93.61524, 93.48286, 93.58395, 93.67625, 93.57587, 93.2342, 91.82615, 
    89.85445, 87.54579, 86.83791, 87.822, 88.24666, 89.31458, 89.74996, 
    90.69863, 91.47652, 91.18156, 89.79252, 84.5489, 75.02878,
  83.29487, 82.3229, 82.08321, 81.38924, 81.28618, 80.38425, 77.33073, 
    72.97006, 70.69319, 70.77297, 71.06277, 71.33669, 72.06532, 73.21803, 
    74.62679, 76.08646, 76.40888, 74.85571, 70.03866, 63.80002,
  74.1011, 74.50536, 74.9297, 74.99176, 74.44745, 73.45003, 72.22772, 
    71.19058, 71.07527, 71.78905, 72.4877, 73.3254, 74.39284, 75.88383, 
    77.39459, 78.26054, 77.08611, 75.78597, 74.36655, 71.85471,
  75.56322, 74.12579, 73.25121, 73.1614, 72.34673, 71.15942, 70.04241, 
    69.40461, 70.21175, 72.00698, 74.6516, 77.60422, 80.107, 81.84768, 
    82.74771, 83.02327, 81.95853, 80.61526, 79.49476, 78.5635,
  76.18433, 74.45004, 72.627, 71.65982, 71.49636, 72.0758, 72.5926, 73.36796, 
    75.61156, 78.7989, 82.20098, 84.86776, 86.81088, 87.96931, 87.8453, 
    86.94646, 85.01112, 82.79234, 81.69091, 80.88367,
  73.16711, 71.77522, 71.28542, 72.66085, 74.73897, 76.60591, 78.18002, 
    79.99298, 82.46709, 85.36757, 87.69522, 89.18459, 89.97424, 90.01562, 
    88.76099, 86.78718, 83.67242, 80.27507, 77.76643, 76.19435,
  71.64504, 74.2802, 77.45116, 79.59138, 80.64577, 81.06041, 79.58099, 
    76.05524, 74.0742, 75.13183, 77.09104, 79.98715, 82.57604, 83.62292, 
    82.884, 81.54295, 77.70529, 72.42114, 68.68298, 67.22098,
  75.75042, 78.52371, 79.8419, 79.07996, 78.1499, 74.44892, 68.18076, 
    64.38321, 63.55277, 62.36189, 61.89007, 63.9155, 67.4728, 70.61604, 
    72.03993, 70.98927, 67.76879, 64.64439, 63.11902, 63.72178,
  73.97388, 74.19803, 73.3336, 72.24086, 72.2293, 68.59734, 66.32502, 
    66.23235, 69.23592, 69.09701, 66.17929, 65.63615, 70.70082, 72.39794, 
    71.46532, 70.58755, 69.46912, 68.17652, 68.04991, 69.59635,
  88.9858, 89.42135, 89.69363, 90.12509, 90.39666, 90.83325, 90.97768, 
    91.36324, 89.9777, 90.45053, 90.79865, 91.14661, 91.36514, 91.64486, 
    92.03632, 92.38174, 91.73917, 91.96878, 92.15668, 92.42601,
  79.16111, 80.49207, 81.93042, 83.45013, 84.8223, 86.29328, 87.6715, 
    88.90804, 85.89934, 87.09655, 88.25091, 89.51325, 90.76306, 91.90435, 
    92.8996, 94.01524, 92.7244, 93.42381, 94.36973, 95.05701,
  77.57041, 79.39301, 81.17284, 83.22619, 85.17868, 87.17082, 89.00359, 
    90.61857, 86.6302, 87.93465, 88.95729, 89.78063, 91.1356, 92.99043, 
    94.57153, 95.70116, 94.658, 95.44688, 96.04865, 96.60079,
  80.38255, 82.71101, 85.06746, 87.32935, 89.51465, 91.38381, 92.80557, 
    93.81648, 91.67931, 92.79682, 93.69231, 94.698, 95.95312, 96.92118, 
    97.54164, 97.7207, 98.35585, 98.27799, 98.20076, 98.02299,
  80.15292, 83.21004, 86.2947, 88.84998, 91.11369, 92.6105, 93.58709, 
    94.64277, 93.64285, 93.84872, 94.39742, 94.64159, 95.49632, 96.38063, 
    97.02287, 97.24178, 99.51064, 99.47217, 99.27309, 98.64761,
  79.3721, 82.63053, 85.24862, 87.29091, 88.47219, 89.23348, 89.78939, 
    90.06762, 85.75269, 85.93648, 86.48732, 87.10805, 87.9828, 89.05282, 
    90.45714, 91.97648, 96.8695, 97.45816, 97.64394, 97.18617,
  92.99684, 91.84456, 91.12887, 91.34769, 91.70437, 92.22652, 91.93797, 
    91.57331, 83.9649, 84.48322, 85.97672, 80.54555, 81.93377, 87.67368, 
    89.25694, 86.96121, 93.4491, 94.59087, 95.63698, 96.00773,
  95.71535, 96.21587, 95.99284, 96.06298, 96.68791, 97.36821, 97.44151, 
    97.4286, 94.83668, 95.056, 95.44305, 92.86206, 93.06783, 95.66938, 
    97.53014, 87.94861, 95.94408, 94.20552, 92.61522, 93.80641,
  94.81257, 94.59109, 94.57195, 94.30253, 93.89073, 94.23661, 93.9318, 
    93.40326, 91.13398, 91.96113, 92.81203, 94.04575, 94.80658, 94.76954, 
    94.41043, 94.54969, 94.58672, 96.71307, 96.72952, 97.22166,
  95.22985, 95.1276, 95.28443, 95.35501, 94.95459, 94.35595, 93.84657, 
    93.4264, 93.18219, 93.33845, 93.65305, 93.81216, 93.72362, 93.56466, 
    93.46323, 93.39062, 93.88409, 94.476, 94.99835, 95.83063,
  95.57659, 95.48354, 95.30968, 94.92601, 94.76143, 94.57787, 94.39719, 
    94.25472, 94.10073, 93.98289, 93.75893, 93.15625, 91.86297, 91.25018, 
    91.66146, 91.86201, 91.68647, 91.94263, 91.69508, 91.83595,
  94.74716, 94.34342, 93.84432, 93.37624, 93.3782, 92.9028, 92.20752, 
    91.32518, 90.18217, 89.42416, 88.76441, 88.00684, 87.5145, 87.94212, 
    88.66488, 90.02771, 89.43056, 89.4821, 87.89331, 84.74616,
  89.69211, 89.06279, 88.6442, 87.96742, 87.42259, 85.69149, 81.54969, 
    77.67605, 75.55907, 75.16994, 74.76401, 74.49462, 75.00536, 76.64954, 
    78.32789, 79.33975, 79.25286, 78.17284, 75.17538, 69.57423,
  78.62371, 78.96103, 79.5337, 79.51805, 78.35289, 76.47487, 74.49378, 
    73.11914, 72.38573, 73.03905, 74.26102, 76.28, 78.83952, 81.40266, 
    83.32326, 83.89005, 82.07729, 80.18026, 78.7432, 76.84431,
  75.93304, 73.79051, 72.73824, 72.53696, 71.82846, 71.18514, 70.5637, 
    70.36122, 70.96055, 73.15816, 76.19108, 79.69289, 82.73113, 84.71862, 
    85.36137, 85.44136, 84.52128, 83.43023, 83.0015, 82.96538,
  71.03696, 69.11665, 67.5106, 67.73072, 68.42247, 69.69874, 70.80616, 
    72.14464, 74.10767, 77.3222, 80.92799, 83.75393, 85.71161, 86.94911, 
    86.84203, 86.29009, 84.88704, 83.10488, 82.61402, 82.30714,
  66.43526, 66.98095, 67.94305, 70.30826, 72.34672, 73.81528, 74.76881, 
    75.79417, 77.01514, 78.89897, 81.07185, 82.95851, 84.17013, 84.84348, 
    84.62616, 83.94448, 81.90811, 79.08051, 76.49001, 74.19189,
  69.55151, 73.17349, 76.41432, 78.83978, 80.04168, 79.93768, 78.80575, 
    75.10007, 70.68539, 70.17944, 71.22581, 72.77467, 74.21042, 75.34959, 
    76.03115, 75.72375, 72.65742, 67.85355, 63.97134, 62.01108,
  76.56474, 78.98997, 79.78302, 79.36734, 79.17807, 76.92293, 71.18398, 
    65.93382, 63.38005, 60.42058, 59.25802, 59.84235, 61.19584, 62.68837, 
    64.26311, 64.58915, 62.72286, 61.14147, 61.83196, 64.02235,
  75.90591, 76.52561, 75.71626, 73.89969, 73.27147, 69.36514, 66.03684, 
    65.02904, 66.40875, 64.41647, 62.02953, 61.01365, 64.98338, 68.55199, 
    69.28062, 69.23628, 68.63747, 69.32966, 72.05657, 75.19295,
  90.89621, 91.11888, 91.36607, 91.64262, 91.93119, 92.20451, 92.45037, 
    92.70847, 91.18864, 91.38273, 91.66953, 91.88114, 92.16753, 92.40924, 
    92.49203, 92.75745, 91.89565, 92.11013, 92.24187, 92.3748,
  84.59005, 85.39179, 86.2606, 87.22884, 88.33301, 89.39272, 90.56348, 
    91.75666, 88.50391, 89.40388, 90.43806, 91.29741, 92.16458, 93.02338, 
    93.77081, 94.56503, 92.63552, 93.2718, 93.8083, 94.1919,
  83.06903, 84.11595, 85.36108, 86.60524, 87.9343, 89.17036, 90.40214, 
    91.67476, 87.47796, 88.84582, 90.08376, 91.08272, 92.19729, 93.18613, 
    94.03543, 94.99174, 93.38298, 94.12642, 95.00422, 95.44625,
  83.87608, 85.68501, 87.54147, 89.14685, 90.54251, 91.92838, 93.33831, 
    94.48409, 91.81031, 92.62904, 93.62047, 94.33203, 95.07731, 95.65137, 
    96.09538, 96.15189, 96.87527, 96.70314, 96.45967, 95.99658,
  83.99622, 86.01778, 88.00352, 88.99454, 90.41269, 91.17407, 92.51815, 
    93.64583, 92.78086, 93.45918, 94.26233, 94.64642, 94.81969, 94.71422, 
    94.88588, 94.99319, 98.59321, 98.44988, 98.12569, 97.1516,
  83.17274, 85.13835, 87.3417, 89.02012, 90.19913, 90.99474, 91.40962, 
    91.48317, 87.12692, 87.04169, 86.66473, 86.69127, 87.2415, 88.25361, 
    89.66856, 90.93256, 97.53595, 97.93425, 97.87296, 97.23208,
  90.66216, 88.69429, 88.11901, 89.17651, 89.90232, 90.49973, 90.67141, 
    89.97643, 81.45244, 81.57899, 80.53134, 79.27445, 80.27641, 84.07332, 
    85.61531, 85.64908, 92.36281, 94.07, 95.41081, 95.96907,
  93.23263, 93.71653, 93.66338, 93.37706, 93.37216, 93.76136, 93.99883, 
    93.70436, 88.55176, 88.71715, 86.08363, 84.26269, 84.94241, 89.61401, 
    91.64219, 79.04579, 90.20477, 92.8325, 92.34267, 93.41473,
  95.14053, 94.99924, 94.88051, 94.84055, 95.06087, 94.74284, 93.94987, 
    93.18885, 91.71724, 91.9664, 92.02541, 90.85475, 89.77107, 89.52118, 
    90.52379, 92.44637, 92.67854, 94.67008, 93.49495, 93.52753,
  96.42583, 96.38694, 96.10419, 95.78692, 95.62304, 95.54242, 95.17258, 
    94.90906, 94.11798, 93.88898, 94.17607, 94.33424, 94.06406, 93.41634, 
    93.05571, 93.56702, 94.8196, 95.7613, 96.34206, 96.53584,
  96.1627, 96.16839, 95.99147, 95.82249, 95.67488, 95.50373, 95.33865, 
    95.01575, 94.52206, 93.77398, 94.04064, 94.58228, 94.85837, 94.51841, 
    94.3875, 94.64278, 94.64363, 94.91036, 95.08933, 95.08098,
  93.93557, 94.42261, 94.58482, 94.58436, 94.89676, 95.09496, 94.99194, 
    94.64466, 93.60168, 93.38242, 93.53943, 93.51518, 93.48721, 93.62813, 
    93.67712, 93.84746, 93.35953, 92.28005, 91.46068, 89.92314,
  88.99575, 89.73719, 90.04398, 90.24363, 90.26369, 89.37785, 86.56447, 
    83.82442, 83.14501, 83.59651, 83.65228, 83.74165, 84.38424, 85.42139, 
    86.03596, 86.27409, 85.34813, 84.17545, 82.57871, 79.18447,
  84.01373, 83.79632, 83.82268, 83.95847, 83.50651, 81.95537, 80.214, 
    78.88189, 78.18343, 78.59587, 79.33303, 80.66345, 82.61027, 84.4487, 
    86.04526, 86.93552, 85.96595, 85.21498, 84.92078, 84.05599,
  80.62612, 77.55188, 76.47598, 76.59835, 75.88335, 74.88898, 74.44121, 
    74.57318, 75.15521, 77.09772, 79.77138, 82.91045, 85.69977, 87.34727, 
    88.03767, 88.30396, 87.69343, 86.76105, 86.71377, 87.21227,
  77.42831, 74.47909, 72.42379, 71.63881, 71.42361, 71.89993, 72.6412, 
    73.78294, 75.65955, 78.83813, 82.21939, 84.95343, 86.72247, 88.13087, 
    88.58691, 88.42464, 87.15964, 85.45715, 85.07806, 85.05977,
  73.09779, 72.00067, 71.8781, 71.95161, 71.83212, 72.27796, 73.40871, 
    75.26768, 76.96142, 78.68926, 80.47295, 82.14854, 83.75208, 85.28403, 
    85.61729, 85.44251, 83.99669, 81.99, 80.56482, 79.75005,
  72.15408, 74.52873, 76.47049, 76.3206, 74.8392, 73.97859, 73.83905, 
    72.1088, 69.16862, 69.22248, 70.73821, 73.13312, 75.6094, 77.1461, 
    78.29886, 78.95924, 76.84203, 72.88489, 70.47279, 70.74837,
  74.53536, 76.49453, 77.11017, 75.95892, 75.07906, 73.39637, 68.9717, 
    63.33126, 59.25502, 57.23076, 56.57352, 58.38041, 61.66562, 64.37842, 
    66.96392, 68.22174, 67.63088, 66.58663, 67.57319, 69.09853,
  72.45463, 71.79242, 70.98843, 70.96592, 71.7412, 68.88503, 64.13661, 
    59.68937, 60.08604, 60.50245, 58.79253, 58.55506, 63.94611, 68.09715, 
    69.61443, 70.03534, 70.37448, 70.31708, 70.44749, 70.81254,
  91.3645, 91.573, 91.67233, 91.89311, 91.97332, 92.19794, 92.36662, 
    92.48856, 91.12385, 91.05939, 91.13206, 91.1679, 91.37714, 91.44641, 
    91.63242, 91.76857, 91.08333, 90.89702, 91.06193, 91.14459,
  85.50427, 86.28353, 86.88442, 87.52236, 88.2956, 89.05345, 89.9842, 
    90.77336, 87.49175, 88.30871, 89.08672, 90.03065, 90.74057, 91.16583, 
    92.06106, 92.69473, 90.71629, 91.15942, 91.40066, 91.91657,
  82.53709, 83.46293, 84.45915, 85.49683, 86.33314, 87.37575, 88.72497, 
    90.05102, 86.10091, 87.43124, 88.33298, 89.07727, 89.92736, 90.76321, 
    91.68478, 92.09344, 90.17944, 90.16369, 90.80061, 90.9724,
  82.57495, 83.90635, 85.08296, 86.1347, 87.24203, 88.37423, 89.38282, 
    90.32861, 87.47168, 88.17715, 88.80773, 89.2641, 89.86105, 90.44386, 
    91.38381, 91.90119, 93.03851, 92.9411, 92.57284, 92.10977,
  81.276, 83.49085, 85.70578, 87.4869, 88.8778, 89.97325, 90.69103, 91.00896, 
    89.16825, 89.62637, 89.67277, 89.55189, 89.66665, 90.04709, 90.28264, 
    90.50839, 95.51801, 95.71612, 94.79672, 93.63401,
  81.24216, 83.61032, 85.90044, 87.8186, 89.09196, 89.69386, 89.81934, 
    89.99222, 85.83409, 85.79588, 85.77153, 86.04309, 86.50374, 87.62961, 
    88.88919, 90.31635, 97.14709, 97.26038, 96.79769, 95.95417,
  85.78819, 84.1634, 84.00113, 84.81228, 85.07527, 85.29876, 85.07829, 
    84.72825, 77.16905, 77.11192, 74.56511, 76.44791, 78.16248, 82.50514, 
    84.92216, 86.20893, 93.78251, 95.95329, 97.01743, 97.19936,
  90.61763, 90.5049, 90.67464, 91.01508, 91.54948, 91.81969, 91.83047, 
    91.57461, 85.73485, 83.8823, 76.97752, 80.17654, 81.30547, 89.16476, 
    86.66296, 79.3889, 79.15128, 92.06599, 91.28747, 93.09615,
  95.33934, 95.09064, 94.46521, 93.60014, 93.13901, 92.32285, 91.07507, 
    89.92318, 86.21002, 85.13565, 84.15936, 83.85056, 84.52587, 86.27717, 
    88.70178, 90.65134, 90.77004, 89.50945, 89.47469, 91.79842,
  96.71568, 96.9405, 96.62625, 96.01116, 94.63091, 93.09302, 91.90439, 
    90.71133, 89.81149, 89.52657, 90.113, 90.99349, 91.4841, 92.04304, 
    93.01663, 93.83064, 93.81626, 94.1026, 94.01377, 93.7495,
  95.81718, 95.5153, 95.64121, 95.47251, 94.99834, 94.53403, 94.1656, 
    93.27493, 92.50094, 91.12013, 90.65867, 90.63244, 90.71528, 90.91431, 
    91.52, 92.35645, 92.9278, 93.30621, 92.90353, 92.75189,
  91.72141, 92.50427, 93.71738, 93.63342, 93.47559, 93.59863, 93.3307, 
    93.14954, 92.88725, 92.23981, 91.39777, 90.81875, 90.46497, 90.33052, 
    90.25976, 90.35394, 90.18944, 89.7117, 88.72306, 87.65096,
  89.50375, 90.91351, 91.7766, 91.89901, 92.01409, 91.40796, 88.97799, 
    86.74698, 86.383, 87.22841, 87.71048, 88.02301, 88.37052, 88.74969, 
    88.98427, 89.32346, 88.90257, 87.8717, 86.0648, 82.07759,
  84.84821, 84.99066, 85.69994, 86.00744, 85.24588, 83.90254, 82.35757, 
    81.21067, 81.24395, 82.03774, 83.08216, 85.12719, 87.26877, 88.88916, 
    90.16446, 90.88161, 89.33301, 87.86965, 86.9704, 85.67596,
  81.54348, 77.96942, 76.12589, 75.82343, 75.48012, 75.54668, 75.99002, 
    76.93822, 78.47679, 80.28609, 82.59045, 85.65743, 88.37455, 89.74089, 
    89.74964, 89.61304, 88.53636, 87.67692, 87.91003, 88.46883,
  76.42992, 73.3195, 71.40477, 71.87323, 73.24374, 75.07585, 77.17126, 
    79.30976, 81.54733, 84.07357, 86.28734, 87.8075, 89.03383, 89.72454, 
    89.27113, 88.75455, 87.88165, 86.98541, 86.99425, 86.57877,
  71.10175, 71.37098, 72.58314, 74.64372, 76.59192, 78.69838, 80.63013, 
    82.08382, 83.64205, 84.84251, 85.80998, 86.66346, 87.53849, 88.58852, 
    88.96047, 88.36542, 86.50208, 84.08064, 82.24412, 80.81959,
  73.02258, 76.3, 78.87653, 79.67557, 79.72928, 80.24851, 79.5901, 77.01684, 
    73.7095, 73.81673, 75.7857, 78.90343, 81.28428, 82.94205, 83.97821, 
    83.59171, 80.63496, 76.14338, 72.83939, 71.29019,
  76.81654, 78.58359, 78.29534, 76.63952, 74.91601, 73.08333, 68.8352, 
    63.99453, 61.63814, 61.30887, 62.42474, 64.58648, 67.72715, 70.201, 
    71.38609, 70.93343, 69.28252, 67.49642, 66.47286, 66.82005,
  72.49437, 71.6625, 69.75641, 68.29561, 68.24616, 67.0891, 65.04065, 
    61.37404, 61.80174, 62.99212, 64.3135, 64.39733, 69.29587, 73.05561, 
    73.36836, 72.57209, 70.97442, 70.47871, 69.79758, 69.53255,
  94.90064, 95.00996, 95.08101, 95.10175, 95.37639, 95.67712, 95.84805, 
    96.23725, 95.14069, 94.37788, 95.10924, 95.12989, 95.1605, 95.26364, 
    95.57732, 95.69822, 95.04958, 94.42651, 95.56937, 95.73177,
  90.06992, 90.67376, 91.58009, 92.28658, 93.00541, 93.41975, 94.09539, 
    94.72912, 91.35695, 92.04633, 92.21258, 92.94515, 93.53311, 94.27477, 
    94.64073, 94.80158, 92.71782, 92.87019, 93.26834, 93.59564,
  86.83752, 87.79669, 89.24849, 90.34772, 91.33627, 92.17843, 93.10141, 
    93.93669, 89.72385, 90.36111, 91.47195, 92.142, 92.7224, 93.39819, 
    93.99378, 94.29298, 92.10622, 92.28614, 92.59753, 92.73886,
  85.21899, 86.60821, 88.54087, 89.64201, 90.42211, 91.08463, 91.90636, 
    92.67364, 89.6377, 90.11754, 91.1161, 91.686, 92.33277, 93.21754, 
    93.67973, 94.12294, 94.7666, 94.44082, 93.62523, 93.06514,
  83.93346, 86.29945, 87.97972, 89.56628, 91.24725, 91.93883, 92.68748, 
    92.86785, 91.13353, 91.66029, 91.88709, 92.385, 92.55491, 92.37224, 
    92.64465, 93.20862, 97.31529, 96.90409, 96.50493, 95.89401,
  82.73397, 85.07328, 86.88776, 88.38313, 89.71446, 90.77895, 91.5893, 
    91.88284, 87.53871, 87.77262, 87.82537, 88.35861, 89.08249, 90.14605, 
    91.13495, 92.41799, 97.86423, 98.00551, 97.74827, 96.93533,
  87.03732, 84.95612, 84.41564, 84.58224, 84.68504, 84.87067, 84.93582, 
    84.90457, 76.95624, 75.83925, 74.41776, 75.65813, 77.24734, 82.23229, 
    85.03012, 86.1011, 93.31994, 95.12951, 96.23892, 96.54712,
  94.18681, 93.97968, 93.37168, 92.64713, 91.51562, 89.43595, 87.19409, 
    84.50672, 74.90685, 71.54491, 70.27235, 76.67512, 77.36029, 80.80839, 
    72.54539, 73.98966, 78.07597, 92.77521, 92.58045, 93.82255,
  95.38631, 94.99299, 94.28216, 93.4137, 92.43939, 90.74946, 88.04623, 
    84.4626, 79.20136, 77.88241, 78.04854, 78.50099, 80.01154, 81.39581, 
    82.2878, 85.9239, 88.51391, 87.66427, 91.04453, 94.43832,
  93.00712, 92.02885, 91.03574, 89.53766, 89.11813, 89.46126, 88.82569, 
    86.94686, 84.65797, 82.71717, 82.64725, 83.14474, 83.76192, 84.41417, 
    84.88572, 85.69563, 86.77204, 87.83794, 88.91284, 89.56184,
  91.16129, 89.79425, 89.28044, 89.09358, 89.34461, 89.94657, 90.30321, 
    89.98326, 88.74429, 87.22488, 86.44852, 86.27288, 86.22276, 85.5984, 
    84.70882, 83.99332, 84.06798, 85.14132, 86.31258, 87.6945,
  92.45391, 92.24512, 92.83517, 92.78235, 92.13048, 91.04652, 89.53388, 
    89.60781, 90.50362, 90.45409, 90.03627, 90.46845, 91.40242, 91.23132, 
    89.3007, 86.85189, 86.13471, 86.26881, 86.26762, 85.78092,
  92.52599, 93.90968, 95.04084, 95.40034, 95.10829, 93.5223, 90.19015, 
    87.53118, 87.19713, 88.26794, 89.06876, 89.69347, 90.67056, 91.68008, 
    91.95544, 91.54601, 90.70938, 89.9871, 89.2302, 86.85352,
  87.8203, 87.88282, 88.32418, 88.40893, 87.72948, 86.52885, 85.29993, 
    84.49593, 84.13013, 84.5996, 85.06063, 85.65453, 87.51411, 90.07048, 
    92.29692, 93.72576, 93.23912, 92.47104, 91.84091, 90.3119,
  84.402, 81.40666, 79.77185, 79.673, 79.49693, 79.69726, 80.29749, 80.93156, 
    81.61623, 82.89632, 84.36444, 85.55179, 87.28263, 89.48326, 91.05511, 
    91.9977, 91.98064, 91.55482, 91.75974, 92.00922,
  79.61, 77.16943, 75.7258, 76.81662, 78.90418, 80.57854, 81.43459, 81.72472, 
    82.22472, 84.39558, 86.68725, 88.13202, 89.40027, 90.35984, 90.78028, 
    90.69949, 90.02717, 89.10295, 89.32232, 88.78273,
  75.10381, 75.1877, 76.32045, 78.80433, 80.22916, 80.42865, 80.50703, 
    80.73585, 80.89033, 82.14877, 83.83013, 85.29885, 85.77946, 86.18816, 
    86.40618, 86.23978, 84.89099, 83.36497, 82.66994, 82.08858,
  77.24128, 78.77406, 79.85229, 79.67782, 78.96619, 78.25731, 77.72816, 
    76.36488, 74.5853, 74.47237, 75.68529, 78.03226, 80.14388, 81.35356, 
    81.68035, 81.38238, 79.24027, 76.50735, 75.27167, 74.97234,
  81.28152, 80.68897, 78.98257, 75.40318, 74.25308, 73.67333, 70.61343, 
    66.79141, 65.3816, 64.5153, 64.99712, 67.80853, 72.35779, 75.00758, 
    76.05123, 75.85421, 74.48849, 72.06738, 70.27673, 70.26532,
  76.79259, 74.37434, 72.11779, 71.18333, 72.29846, 71.74786, 68.35709, 
    61.58953, 62.47335, 64.20592, 64.88162, 66.53403, 71.55174, 75.10848, 
    75.22465, 75.17352, 74.2563, 72.58195, 72.41462, 74.92426,
  93.216, 93.51062, 93.789, 94.06239, 94.49396, 94.75712, 94.92636, 95.15638, 
    93.63091, 94.13532, 94.17456, 94.34935, 94.94543, 95.17426, 95.51659, 
    94.87414, 95.4415, 94.61515, 94.97452, 95.00442,
  88.97779, 89.85695, 90.7765, 91.64599, 92.56039, 93.47754, 94.23036, 
    94.94672, 91.4035, 92.06362, 92.74107, 93.40923, 94.22253, 94.9411, 
    95.70839, 96.22915, 94.13529, 94.80077, 95.50822, 96.22432,
  84.75642, 86.35967, 88.12784, 89.93417, 91.53645, 93.13905, 94.53223, 
    95.56105, 91.2412, 92.1717, 92.96066, 93.85765, 94.69868, 95.44509, 
    96.15118, 96.82774, 95.03838, 95.75444, 96.42094, 96.93476,
  86.43343, 88.34901, 90.12505, 91.71494, 93.11809, 94.30839, 95.48973, 
    96.61714, 94.33985, 94.83659, 95.46133, 95.95019, 96.52157, 96.89012, 
    97.13544, 97.31297, 98.01559, 98.08018, 98.06102, 97.97695,
  86.11224, 88.21268, 90.27713, 92.4492, 94.19518, 95.34867, 96.23286, 
    96.88295, 95.99525, 96.51287, 96.9637, 97.10341, 97.1278, 96.78065, 
    96.51015, 96.26449, 98.87968, 98.53809, 98.12453, 97.46763,
  87.2118, 89.41763, 91.59333, 92.87872, 94.01726, 94.94121, 95.30289, 
    95.65471, 91.05128, 90.87875, 90.8238, 91.25923, 91.53782, 91.82629, 
    92.32576, 92.69979, 97.90283, 97.502, 96.62711, 95.30042,
  93.80304, 92.21922, 91.83633, 92.02191, 90.29782, 89.62868, 88.62254, 
    88.16432, 80.39298, 79.97565, 79.87415, 82.18704, 83.87831, 88.09332, 
    90.73753, 89.74113, 94.65026, 95.03704, 95.09872, 94.96138,
  80.47141, 77.70677, 75.26943, 74.4869, 71.48505, 69.94061, 68.27101, 
    67.26982, 61.52334, 60.16146, 59.71165, 68.15359, 75.03677, 83.55528, 
    82.05031, 85.07533, 89.34256, 91.21207, 89.10944, 88.75771,
  74.61462, 74.50706, 74.19028, 73.69572, 73.32972, 73.18715, 72.50208, 
    71.6451, 69.33759, 70.59086, 72.48738, 74.7306, 77.92234, 82.49602, 
    84.78788, 85.48773, 83.64599, 82.44233, 87.6806, 90.92067,
  77.30231, 77.07834, 76.95487, 77.0026, 77.69582, 78.30352, 78.32803, 
    77.55229, 76.34258, 76.25141, 77.94728, 80.45915, 82.89703, 85.08298, 
    86.95464, 88.41443, 90.0218, 90.9558, 90.85185, 90.60954,
  81.65134, 80.84237, 80.71913, 80.6349, 81.15538, 81.94046, 82.00108, 
    81.44781, 80.82392, 80.43937, 81.34074, 83.4417, 85.42754, 86.81457, 
    87.85324, 88.2562, 89.22237, 90.34833, 91.16629, 91.92946,
  83.37442, 83.02296, 83.56842, 84.46716, 85.29488, 84.60869, 83.18311, 
    82.24489, 83.38145, 84.72242, 85.57249, 87.24186, 89.15244, 91.08679, 
    91.86066, 90.93749, 91.32639, 91.69442, 91.12396, 90.18413,
  86.65727, 87.35411, 87.56695, 87.79165, 87.72646, 86.00437, 82.8539, 
    81.17216, 82.75083, 85.71791, 88.09158, 90.16562, 91.9088, 93.29776, 
    94.32468, 94.97968, 94.87518, 93.87952, 92.48331, 89.96156,
  84.26029, 83.56408, 82.87572, 81.53337, 79.9878, 78.7864, 78.37675, 
    79.42032, 82.78922, 85.88817, 88.03411, 90.01813, 91.63015, 93.01389, 
    94.53947, 95.75605, 95.62463, 94.9347, 94.11761, 92.69372,
  80.01603, 76.53326, 74.40072, 73.62858, 73.07848, 73.72451, 75.76421, 
    78.48583, 81.81818, 84.33157, 86.83963, 89.46043, 91.11459, 92.52654, 
    93.97279, 94.7067, 94.77562, 94.58833, 94.86826, 94.88205,
  74.72959, 71.53463, 69.83343, 70.49773, 72.2342, 74.67789, 77.42339, 
    79.48242, 81.78035, 84.55872, 86.98445, 88.86532, 90.41975, 92.11609, 
    93.21838, 93.69218, 93.42017, 92.93401, 93.35341, 93.08413,
  70.7744, 70.41328, 70.83951, 72.41956, 74.5713, 76.30545, 76.848, 77.01794, 
    78.50288, 81.17908, 83.24457, 84.77047, 86.7328, 88.59637, 89.21707, 
    88.86608, 87.60991, 86.15279, 85.97172, 86.51274,
  73.10735, 74.77612, 75.4995, 75.53365, 75.23713, 74.12589, 72.23372, 
    69.49979, 68.92664, 70.48698, 73.06438, 76.41516, 79.70693, 82.06184, 
    82.52037, 82.0518, 80.15067, 77.72237, 76.35593, 77.33678,
  74.43034, 75.54536, 74.61425, 72.07451, 69.95, 67.35821, 62.92334, 
    60.43759, 61.25076, 61.84196, 63.81509, 67.1236, 70.85104, 73.39632, 
    73.94308, 72.70277, 71.5181, 70.84182, 71.33753, 72.15327,
  67.95904, 67.16582, 65.37699, 63.93146, 64.54757, 63.46764, 62.78434, 
    61.99448, 64.4307, 65.90632, 67.31347, 68.69995, 72.029, 74.06059, 
    72.63055, 71.04193, 70.74175, 71.39549, 72.40318, 73.34933,
  89.79278, 90.37881, 90.84624, 91.28751, 91.77792, 92.19527, 92.77354, 
    93.0704, 91.79471, 91.96838, 92.46144, 92.72598, 93.05687, 93.37714, 
    93.72061, 93.89969, 93.34924, 93.33206, 93.54109, 93.43903,
  84.50379, 85.82011, 87.03454, 88.21743, 89.26495, 90.21261, 91.00681, 
    91.74123, 88.44184, 89.12884, 89.64782, 90.06282, 90.8521, 91.84962, 
    92.94142, 94.03995, 92.40247, 93.15495, 94.60784, 95.7111,
  84.81741, 86.48399, 88.21575, 89.75912, 91.17986, 92.26382, 93.08364, 
    93.60173, 89.21716, 89.84933, 90.38229, 91.88002, 92.8958, 94.03183, 
    95.06798, 95.8733, 95.17502, 96.08081, 97.08924, 97.80367,
  83.2972, 85.15878, 86.99529, 88.72662, 90.19515, 91.55212, 92.52174, 
    93.40816, 91.23263, 92.54955, 92.90449, 94.27661, 95.17411, 96.13899, 
    97.44017, 97.91475, 98.08382, 98.25446, 98.50152, 98.30161,
  79.12604, 81.11093, 82.88255, 84.84923, 86.59763, 88.19781, 89.28374, 
    90.96352, 90.91696, 92.57832, 93.83304, 94.96735, 95.84206, 96.28783, 
    96.55592, 95.97031, 97.71371, 97.96048, 98.0106, 97.53111,
  79.57648, 82.00039, 84.00725, 85.42104, 86.2607, 87.08006, 87.94465, 
    88.69449, 84.92491, 85.3433, 85.76184, 86.6475, 87.4003, 87.97797, 
    88.51122, 89.48006, 95.42224, 96.08701, 95.60403, 95.38906,
  89.24516, 88.11227, 88.20884, 88.64435, 88.93238, 90.60493, 90.37812, 
    90.32917, 82.90945, 82.65495, 83.66127, 78.01855, 79.41806, 84.52693, 
    87.54865, 84.1693, 89.94269, 91.32874, 92.20176, 93.17925,
  79.57878, 76.01755, 73.61486, 69.80401, 68.45731, 70.54015, 69.81189, 
    68.76951, 62.58468, 62.07023, 67.53337, 75.5619, 78.69382, 85.45087, 
    89.5711, 91.34069, 93.37431, 91.59051, 88.89849, 88.21432,
  70.53488, 70.5442, 69.98475, 69.05635, 68.50446, 68.9865, 70.45495, 
    72.35147, 71.58754, 72.11631, 71.91898, 71.38208, 72.82343, 76.47874, 
    79.76989, 82.03355, 84.82838, 87.51237, 89.01825, 90.35078,
  77.11404, 77.42894, 77.48676, 77.47517, 77.47393, 77.77013, 78.27209, 
    78.4098, 79.19626, 79.87354, 80.02749, 80.07943, 80.22679, 80.71193, 
    81.29959, 81.69061, 81.49001, 81.17103, 80.99521, 80.39266,
  80.91624, 81.44832, 81.93004, 82.20585, 82.51162, 82.47764, 82.6323, 
    82.83749, 83.24744, 83.46022, 83.96711, 84.756, 85.22659, 85.68216, 
    85.90187, 86.10682, 85.60508, 84.97642, 84.51593, 84.26587,
  83.26441, 83.80345, 84.60149, 85.31387, 85.68062, 84.62566, 83.15912, 
    83.47244, 85.57837, 87.10149, 87.68399, 88.06184, 88.60851, 88.99815, 
    89.11066, 89.01093, 87.98843, 86.96763, 85.19171, 83.5013,
  83.6033, 84.98266, 85.67326, 86.11816, 86.14242, 85.08582, 83.06745, 
    81.8462, 82.80471, 84.23855, 85.48976, 86.77442, 88.04292, 89.07376, 
    89.94546, 90.66969, 89.5727, 88.00218, 86.16892, 83.53802,
  80.96968, 80.56503, 80.55604, 80.78481, 80.4938, 79.89896, 79.33892, 
    79.28604, 80.08965, 81.41226, 83.10455, 84.85847, 86.3838, 87.48335, 
    88.54082, 89.06028, 87.84209, 87.04095, 86.55164, 85.18182,
  79.63506, 76.71326, 75.408, 75.67774, 75.75038, 75.85552, 76.23798, 
    77.35287, 79.49377, 81.63569, 83.4757, 85.22535, 86.66631, 87.26272, 
    87.27354, 87.03976, 85.56626, 84.42129, 84.65079, 84.91421,
  76.31187, 73.80573, 72.69727, 74.20355, 76.02271, 77.61665, 79.28822, 
    81.07729, 82.61541, 83.604, 84.5099, 85.67027, 86.78809, 87.00987, 
    86.27365, 85.70525, 84.02746, 82.27774, 81.97807, 80.64091,
  73.60911, 74.41924, 76.30058, 78.76736, 80.02112, 80.73661, 81.27076, 
    81.40185, 82.25658, 83.27487, 84.01122, 84.50988, 84.81628, 84.64581, 
    84.69954, 84.02905, 81.93338, 79.19004, 76.83179, 74.68038,
  77.52993, 79.7002, 81.22529, 81.35121, 79.95695, 78.85426, 78.45315, 
    77.15611, 76.445, 76.98684, 77.92998, 79.55824, 80.84178, 80.8673, 
    80.33311, 79.17357, 76.91196, 74.05534, 72.26131, 71.33239,
  77.96581, 78.47338, 77.26288, 75.13734, 74.27358, 74.13857, 72.48808, 
    70.31044, 69.37407, 67.96851, 66.61884, 66.50686, 67.63235, 68.59193, 
    69.91575, 70.76519, 71.42197, 71.62648, 72.31139, 71.75679,
  69.56062, 68.38315, 66.82086, 66.78863, 69.19053, 71.48899, 72.40832, 
    68.80007, 68.6744, 68.15332, 65.68047, 63.85214, 66.10426, 70.65089, 
    73.27699, 73.83241, 73.80519, 73.56245, 73.74154, 72.96153,
  92.1509, 92.47922, 92.78604, 92.9416, 93.43333, 93.36813, 93.94291, 
    93.94337, 92.66093, 92.89922, 93.17401, 93.62741, 94.06394, 94.42846, 
    94.6459, 95.28361, 94.26261, 94.74635, 94.67545, 95.32315,
  86.34003, 87.73792, 89.0783, 90.67628, 92.27706, 93.94343, 94.88348, 
    95.61666, 92.29687, 93.34605, 94.05518, 94.36356, 94.95261, 95.49216, 
    96.29266, 96.86999, 95.52209, 96.22078, 96.9508, 97.48348,
  88.46748, 90.49299, 92.44296, 93.86613, 94.80479, 95.44716, 95.99785, 
    96.32353, 91.85777, 93.16527, 94.87513, 96.27115, 97.00442, 97.64667, 
    98.22755, 98.39138, 97.55653, 97.8643, 98.12475, 98.24935,
  87.58758, 90.06383, 91.96062, 93.86033, 94.99348, 95.96637, 96.78468, 
    97.263, 95.87243, 97.05312, 97.95033, 98.74782, 99.16679, 99.46056, 
    99.42163, 99.74187, 99.97818, 99.96271, 99.75571, 99.30542,
  86.02782, 89.10584, 91.71903, 93.69155, 94.84707, 95.27446, 95.40157, 
    94.01119, 92.69804, 92.51897, 93.21578, 94.28227, 95.38741, 96.24226, 
    96.77219, 97.15907, 98.96427, 99.07253, 98.61249, 98.28286,
  86.85065, 89.6467, 91.89108, 92.74184, 92.7908, 92.22177, 91.09188, 
    90.01849, 85.78457, 85.99502, 86.73858, 87.63344, 88.35235, 89.42884, 
    90.31464, 90.96222, 96.58284, 97.33385, 97.92881, 97.55293,
  97.70763, 96.47759, 96.38071, 95.79133, 94.64653, 94.07471, 93.31896, 
    92.3814, 85.18241, 85.57598, 87.38814, 79.25886, 80.30389, 86.47298, 
    89.15688, 85.35068, 91.36413, 93.18764, 94.53224, 95.4276,
  95.21188, 94.57956, 93.08287, 91.05466, 89.1101, 87.96649, 88.19984, 
    89.42628, 84.16132, 86.36071, 90.00322, 87.67043, 88.6624, 92.56511, 
    93.82767, 95.56513, 95.39212, 95.16305, 92.65701, 93.79205,
  70.77306, 68.36935, 67.67353, 67.32683, 67.81615, 69.00539, 68.97746, 
    68.04552, 65.08203, 67.17127, 70.86951, 77.58215, 84.66106, 90.55525, 
    93.03986, 95.39828, 96.79596, 97.8955, 98.34296, 98.24023,
  69.1435, 69.96334, 71.27856, 72.15461, 72.97527, 73.65043, 73.81712, 
    73.15318, 71.76665, 70.50961, 69.97007, 70.38229, 71.72931, 74.24483, 
    75.52213, 75.5317, 76.51327, 77.82415, 80.41833, 84.27782,
  74.1205, 75.02709, 76.01174, 76.76492, 77.33358, 77.6422, 78.07654, 
    78.34727, 78.11507, 77.29336, 76.80334, 76.92184, 77.47813, 77.95372, 
    78.21468, 78.22069, 77.69842, 76.79279, 76.58381, 77.11197,
  79.77225, 80.25014, 80.38916, 80.29462, 80.2532, 78.67474, 77.46124, 
    78.25684, 80.61267, 82.04851, 82.25126, 82.29808, 82.88591, 83.70813, 
    84.13673, 83.95316, 83.17665, 81.75345, 79.79922, 78.26664,
  80.67493, 81.87469, 82.48022, 82.48722, 82.28519, 81.00954, 78.53385, 
    76.87337, 77.2622, 78.52731, 79.93253, 81.30635, 82.97153, 85.07201, 
    86.94083, 87.85825, 87.75938, 86.45996, 84.59982, 81.69284,
  76.73793, 76.77984, 77.01991, 77.0884, 76.54785, 75.57635, 74.4838, 
    73.82414, 74.53901, 76.11497, 78.20918, 80.92307, 84.00097, 86.86723, 
    89.40571, 90.8242, 90.19323, 89.0823, 88.20142, 86.73849,
  77.09907, 74.17075, 72.19415, 71.52142, 70.75912, 70.3239, 70.30522, 
    70.91906, 73.36388, 76.381, 79.81072, 83.21574, 85.84622, 87.66133, 
    88.7943, 89.33173, 88.25683, 86.96069, 87.14232, 87.50299,
  74.41276, 70.64822, 67.84197, 68.0872, 69.67619, 71.16582, 72.38897, 
    74.55772, 78.27148, 81.4499, 83.95437, 85.90337, 87.21224, 87.84589, 
    87.81939, 87.5956, 86.50665, 85.55251, 86.18161, 85.96653,
  68.00421, 67.53833, 69.01143, 72.1477, 74.56783, 75.7681, 76.35052, 
    76.98061, 78.80279, 81.17322, 82.79155, 83.85787, 84.75467, 84.95809, 
    84.88222, 85.01089, 83.90862, 82.07978, 80.84544, 80.4499,
  68.5594, 70.96941, 73.58348, 74.86653, 74.35104, 72.97656, 70.42741, 
    67.06526, 64.81364, 66.47118, 70.37269, 75.03369, 79.06978, 81.1698, 
    82.37658, 82.12482, 79.65471, 75.57366, 73.69397, 73.98529,
  69.96117, 71.05347, 70.67908, 68.9779, 66.82713, 64.05182, 60.13258, 
    58.04848, 58.20843, 58.24718, 60.28251, 65.31539, 71.64214, 75.16063, 
    76.21164, 75.0595, 72.76579, 70.9439, 70.9183, 71.995,
  65.06496, 63.26559, 61.37787, 61.4031, 62.98011, 62.32104, 63.36922, 
    64.05184, 65.36583, 66.78902, 65.16712, 67.2127, 73.8317, 77.30964, 
    75.76283, 73.57456, 71.80347, 70.99984, 72.19592, 73.15749,
  92.73816, 93.36729, 93.69086, 94.06555, 94.31395, 94.65488, 95.00951, 
    95.32661, 93.87023, 94.33353, 94.70605, 95.01334, 95.28855, 95.63437, 
    96.02279, 96.13508, 95.37886, 95.75971, 95.93408, 95.97202,
  88.33485, 89.41888, 90.16246, 91.23414, 92.19819, 93.22892, 94.20995, 
    95.2645, 91.84321, 92.71059, 93.3244, 94.51392, 95.46542, 96.02596, 
    96.54281, 97.13706, 95.82472, 96.32922, 96.67727, 97.25043,
  86.27853, 87.75147, 89.20423, 90.62852, 91.86864, 92.94179, 93.75928, 
    94.61077, 90.27551, 91.79277, 93.17421, 94.43695, 94.96367, 95.35143, 
    95.87926, 96.3242, 95.67129, 96.05199, 96.80483, 97.04345,
  85.6271, 87.28356, 88.91502, 90.38824, 91.85424, 93.27074, 94.0119, 
    94.49979, 92.13921, 93.03149, 94.3899, 95.80059, 97.1008, 98.24787, 
    98.8688, 99.07267, 99.04839, 98.72356, 98.1918, 97.05173,
  80.79221, 82.73937, 84.94617, 86.26524, 86.90136, 87.34753, 87.46362, 
    87.39724, 86.96584, 87.94042, 89.51961, 91.5353, 92.87983, 94.72472, 
    96.7474, 97.57063, 99.02068, 98.97736, 98.97268, 99.01024,
  78.61961, 81.04375, 83.10923, 84.66141, 85.35304, 85.46783, 85.41589, 
    84.60178, 80.77804, 81.36826, 82.46901, 83.87864, 85.25755, 86.52981, 
    87.86353, 89.646, 96.9424, 97.83731, 97.8329, 97.35823,
  92.55454, 88.13053, 87.40472, 87.23586, 87.37325, 88.16345, 87.82537, 
    86.63633, 78.3765, 77.36389, 78.81843, 74.26379, 75.31277, 79.16395, 
    82.3456, 80.82821, 87.14478, 89.362, 91.15587, 92.05394,
  97.55847, 96.48278, 95.08381, 94.37318, 94.39957, 95.00018, 95.09574, 
    94.69508, 88.12479, 88.23335, 91.04628, 83.75058, 82.39282, 86.16633, 
    91.7859, 92.98334, 93.56952, 91.76167, 89.36505, 90.49986,
  95.12081, 93.41819, 90.50536, 88.97348, 88.01745, 88.32037, 88.6853, 
    89.73515, 89.88182, 93.10722, 94.76971, 95.58704, 95.48777, 94.89742, 
    93.92292, 93.63776, 94.88767, 96.56228, 97.55199, 97.14877,
  86.81734, 83.387, 78.80066, 75.69331, 74.22327, 72.21415, 70.25212, 
    72.67347, 76.38604, 78.36546, 81.37916, 86.36495, 89.13102, 90.57348, 
    90.42374, 89.73675, 89.11744, 89.89061, 92.16722, 94.59732,
  77.95338, 78.4802, 77.46521, 75.77059, 72.74072, 69.46677, 68.61296, 
    68.99946, 69.89797, 71.06297, 72.88248, 75.10216, 77.27509, 78.47164, 
    78.20525, 77.36568, 76.13506, 74.52143, 73.48296, 74.02187,
  74.27925, 74.5815, 74.25751, 73.4048, 72.89632, 71.51342, 70.13556, 
    70.59162, 72.30955, 74.60228, 76.3214, 77.72585, 78.9071, 80.21107, 
    80.91865, 80.51354, 79.60463, 77.94645, 75.71638, 73.83804,
  76.68177, 76.98859, 76.74562, 76.0527, 75.44585, 74.40178, 72.74075, 
    71.70972, 71.7287, 73.13723, 74.71301, 76.04753, 76.85675, 78.11281, 
    79.72974, 80.95178, 81.21, 80.41427, 79.29321, 77.54282,
  76.79292, 76.18129, 75.62177, 74.88414, 73.6885, 72.21393, 70.71922, 
    69.84589, 69.11095, 69.14598, 69.99841, 71.57238, 73.63079, 75.95487, 
    78.76269, 81.12345, 81.71196, 81.48155, 81.29144, 80.12431,
  77.15519, 74.28594, 71.7895, 70.1809, 68.58612, 66.7775, 65.56381, 
    65.06843, 65.67664, 67.61377, 70.70541, 74.13699, 77.41574, 80.10669, 
    82.23109, 83.39069, 82.95945, 81.78255, 82.11047, 82.86398,
  74.24647, 70.69541, 66.83629, 65.29087, 65.71995, 66.55448, 67.35001, 
    68.71671, 72.17323, 76.10339, 79.7743, 82.87244, 85.14935, 86.22394, 
    85.90228, 84.94044, 83.41151, 82.07088, 83.18419, 83.49007,
  69.48212, 68.58279, 69.35592, 71.24619, 72.88068, 74.06171, 75.01589, 
    76.08937, 77.94293, 80.75832, 82.61286, 83.39157, 83.80418, 84.20815, 
    83.71519, 82.83701, 81.35932, 79.52287, 78.69299, 78.6115,
  71.1186, 74.23594, 77.50877, 78.72762, 77.99516, 76.84792, 73.89217, 
    69.60857, 67.45979, 68.47183, 70.10012, 72.33989, 74.15619, 75.59614, 
    76.79097, 77.45808, 76.23511, 74.09062, 73.04171, 72.88757,
  73.58972, 75.84557, 76.55463, 76.23659, 74.9563, 70.21186, 63.47978, 
    59.43633, 58.04411, 56.39864, 55.3165, 56.6959, 59.96147, 63.88914, 
    67.84066, 69.88289, 70.94794, 71.60458, 72.47061, 73.16376,
  69.78126, 68.65292, 67.50025, 67.92507, 68.67879, 65.60644, 64.74046, 
    65.43841, 65.28607, 63.72516, 57.12598, 57.20245, 63.43385, 69.08446, 
    71.66192, 73.20412, 73.98795, 74.53982, 75.17136, 74.27499,
  90.89503, 91.32497, 91.60706, 91.80373, 92.02844, 92.10624, 92.59859, 
    92.93288, 91.66312, 92.18697, 92.54333, 92.97706, 93.37431, 93.87121, 
    94.26491, 94.57002, 93.88563, 94.26356, 94.57425, 94.72278,
  87.32605, 88.25643, 89.10403, 90.00215, 91.06298, 92.21971, 93.46282, 
    94.65732, 91.64652, 92.56804, 93.68418, 94.44693, 95.08447, 95.46259, 
    95.7707, 96.22617, 94.7532, 95.42282, 96.05388, 96.43637,
  88.23593, 89.56976, 90.67647, 91.37772, 92.28933, 93.36485, 94.49519, 
    95.64948, 91.9231, 92.66587, 93.51585, 94.58913, 95.8687, 95.51612, 
    95.55891, 96.30222, 96.14368, 97.13409, 97.69924, 98.40812,
  87.50043, 89.93722, 92.24789, 93.87999, 94.86498, 95.76873, 96.38215, 
    96.79099, 95.1395, 95.27818, 95.39866, 94.77626, 94.82367, 95.30645, 
    95.96176, 97.17538, 98.49734, 99.3025, 98.67153, 97.39704,
  82.25327, 83.88755, 85.99963, 88.65113, 91.33241, 92.72771, 93.14926, 
    93.16695, 92.78705, 92.88011, 92.35917, 91.91406, 92.14445, 93.15054, 
    94.02398, 95.11514, 97.88181, 98.41503, 98.76497, 97.85664,
  80.00447, 81.81201, 83.27109, 84.97996, 86.5563, 87.61384, 87.76379, 
    87.4778, 84.17276, 85.31038, 86.32766, 87.54256, 89.02065, 90.77468, 
    92.04317, 93.17491, 98.14297, 98.28336, 98.04768, 97.1527,
  93.36369, 88.33085, 89.27205, 90.11233, 90.22041, 90.09583, 89.44617, 
    89.48206, 81.81346, 83.07912, 86.07246, 81.80209, 83.9008, 89.45882, 
    91.29783, 90.67464, 95.25126, 96.36842, 96.62243, 95.79838,
  97.31618, 96.88737, 96.49032, 95.84528, 95.51518, 94.78066, 94.4207, 
    94.63351, 91.55205, 93.67634, 95.83462, 93.1638, 93.39223, 94.87704, 
    95.30847, 96.48363, 96.37218, 97.79091, 93.70528, 94.87538,
  94.65803, 94.7355, 94.5396, 94.58878, 95.08025, 95.49854, 95.51878, 
    95.16917, 94.40589, 95.74131, 97.49903, 98.17392, 97.80018, 97.35585, 
    97.67538, 97.87263, 98.84584, 99.2644, 99.13718, 98.76852,
  95.13779, 94.46685, 94.89259, 95.58025, 96.10058, 95.89204, 95.09522, 
    95.30145, 95.41898, 95.78387, 96.61171, 97.51837, 97.17725, 96.68285, 
    96.59712, 96.78488, 97.4461, 97.98081, 98.01367, 98.15735,
  96.06234, 96.69871, 96.69679, 96.21033, 95.43707, 91.02518, 85.59448, 
    84.11619, 85.0415, 87.40789, 89.61104, 90.68695, 90.81075, 90.09887, 
    88.69179, 85.58904, 80.8801, 75.18356, 72.66969, 74.15569,
  82.94685, 85.39324, 86.71391, 85.78831, 83.3244, 78.33805, 75.19891, 
    75.07453, 76.64102, 77.76324, 78.13994, 78.04797, 78.01006, 78.4111, 
    78.15598, 76.7688, 75.45522, 74.13692, 72.41009, 71.08441,
  84.32378, 85.0472, 85.52727, 85.64379, 85.35844, 83.48572, 80.97904, 
    79.44211, 79.88431, 80.8531, 81.34691, 81.89549, 82.57151, 83.31696, 
    84.00407, 84.26267, 83.12421, 81.36955, 79.5685, 76.74966,
  81.84706, 81.1494, 81.10867, 82.03483, 82.31668, 81.80685, 81.08517, 
    80.94548, 81.60521, 82.12109, 82.29322, 82.87508, 84.25862, 85.95235, 
    87.55974, 88.60015, 87.1319, 85.50407, 84.14862, 82.0746,
  77.75754, 74.44892, 72.94573, 73.47004, 73.34033, 73.54954, 74.29119, 
    75.83276, 78.30373, 80.26862, 82.32596, 84.78226, 86.84216, 88.31464, 
    88.84268, 88.63891, 86.96043, 84.88219, 83.6146, 83.03252,
  72.19866, 68.52728, 65.07634, 64.48803, 65.74221, 68.39807, 71.4249, 
    74.8688, 79.56214, 83.51044, 86.73906, 88.94471, 90.20382, 90.50188, 
    89.04313, 86.78384, 83.55717, 81.09429, 81.0115, 80.74593,
  63.51044, 61.77928, 62.99557, 67.13269, 71.06809, 74.67593, 77.89478, 
    81.0156, 84.819, 87.56899, 89.06564, 89.6584, 89.88209, 89.63016, 
    88.14736, 85.60944, 82.0719, 79.21498, 77.43362, 76.00394,
  64.15341, 68.05822, 72.84027, 76.89373, 79.09299, 80.26793, 78.74328, 
    75.60494, 74.42358, 75.82304, 78.18442, 80.86199, 82.90429, 83.22869, 
    82.6655, 81.17861, 77.46443, 72.90141, 70.08612, 68.99479,
  71.99527, 75.08354, 76.79375, 77.57905, 77.60799, 73.26781, 66.25611, 
    62.07297, 61.09129, 59.08176, 58.35947, 60.24057, 63.90074, 66.95718, 
    67.66525, 67.1248, 66.31834, 66.20871, 67.30427, 68.73232,
  69.93742, 69.7103, 69.27615, 70.42594, 71.30301, 67.35316, 65.96633, 
    66.122, 66.91823, 64.31965, 57.35582, 57.16715, 62.2882, 66.18121, 
    66.57986, 66.81626, 68.40799, 70.02795, 71.12891, 70.9048,
  91.86416, 91.94788, 92.35681, 92.46732, 92.71998, 93.12737, 93.28974, 
    93.62265, 92.26591, 92.64647, 93.01614, 93.20046, 93.64958, 94.09109, 
    94.64189, 94.93652, 94.38986, 94.60286, 94.66582, 94.94074,
  86.43339, 87.86991, 89.13162, 90.3647, 91.39756, 92.28436, 93.19794, 
    93.82683, 90.1469, 90.9369, 91.76517, 92.47111, 92.96478, 93.32269, 
    93.72425, 94.2217, 93.22806, 94.19464, 96.21848, 96.95283,
  91.52789, 92.51314, 93.35435, 94.11354, 94.63834, 94.86472, 95.12748, 
    95.27946, 90.80096, 91.61617, 92.46821, 93.59792, 95.32163, 96.76898, 
    97.70712, 98.06458, 97.24444, 97.66802, 98.02302, 98.57449,
  89.32896, 91.50015, 92.93855, 94.07615, 94.87164, 95.62183, 96.3949, 
    96.67976, 95.36484, 96.4229, 96.92516, 97.37255, 97.83807, 98.17416, 
    98.60964, 98.7988, 98.99178, 98.96655, 98.60967, 97.84619,
  87.58652, 90.21882, 92.45762, 93.52962, 92.92955, 93.14032, 93.38831, 
    93.3425, 92.02536, 91.86536, 92.45219, 93.17215, 94.04031, 95.13493, 
    96.38865, 97.35342, 98.2386, 97.943, 97.46552, 97.37858,
  83.17204, 85.08608, 86.99761, 88.31211, 88.47733, 87.96884, 87.94267, 
    87.8537, 83.58051, 84.25444, 85.18191, 86.16354, 87.40843, 88.43565, 
    88.93314, 89.43366, 95.78157, 96.86234, 97.42853, 97.28535,
  94.40118, 92.01391, 91.69241, 91.10684, 88.96226, 87.57042, 86.99899, 
    86.14531, 78.07439, 78.87917, 80.85889, 75.93344, 77.19537, 82.13329, 
    83.73523, 81.84191, 86.87659, 88.2085, 89.42658, 89.89413,
  98.1888, 97.24693, 96.24709, 95.08498, 93.90452, 93.86198, 93.33721, 
    92.85464, 88.84218, 90.96706, 92.91846, 89.13174, 87.57891, 89.67891, 
    91.44029, 90.4044, 91.43131, 87.69032, 86.67567, 87.42791,
  98.33624, 98.45329, 98.68967, 98.51659, 98.20242, 98.14562, 97.59196, 
    96.60587, 93.92171, 93.70004, 94.55052, 95.97034, 96.41224, 96.7823, 
    96.94202, 97.12149, 97.50748, 98.01557, 97.11319, 95.81797,
  97.67355, 98.01227, 98.19881, 98.28868, 98.46585, 97.92423, 97.13302, 
    96.17395, 96.81867, 96.95219, 97.18034, 97.80849, 98.41897, 98.3849, 
    98.46392, 98.48859, 98.31151, 98.24268, 97.9661, 98.07344,
  97.52465, 97.52612, 97.2466, 96.98891, 96.92647, 94.93573, 92.12641, 
    92.75719, 95.01813, 95.98525, 96.23454, 96.66383, 97.07315, 97.41154, 
    97.79855, 97.83215, 97.21226, 93.52736, 81.43838, 75.15238,
  90.6338, 91.89018, 92.11729, 91.444, 88.21819, 76.44162, 67.00648, 
    66.68871, 71.03253, 74.17288, 74.99246, 75.23645, 76.35431, 78.44244, 
    82.25446, 84.6329, 82.68224, 71.92828, 61.99562, 58.16951,
  70.67503, 72.02916, 71.9438, 71.50063, 71.41319, 69.98882, 68.16038, 
    67.10169, 67.23257, 68.48618, 69.66795, 70.44179, 71.19587, 72.16382, 
    73.37697, 74.77729, 74.14881, 72.23713, 70.15369, 67.73012,
  65.77337, 64.83869, 64.61319, 65.34972, 65.81952, 65.53623, 64.89703, 
    64.51677, 65.37115, 67.55559, 69.55792, 71.63375, 73.83518, 76.44501, 
    79.25848, 81.39967, 80.98322, 80.42446, 80.00324, 78.61655,
  65.32689, 61.64551, 59.35399, 59.31601, 58.83395, 58.06224, 57.88971, 
    58.6496, 60.91548, 63.95967, 67.60534, 71.89213, 76.17168, 79.96299, 
    82.55604, 83.85214, 83.22751, 82.10689, 81.65544, 81.87231,
  62.73829, 58.31649, 54.59621, 53.67055, 53.92221, 55.05518, 57.03729, 
    59.30372, 62.81891, 67.36767, 72.54729, 77.42435, 81.28154, 84.43453, 
    86.00908, 85.45322, 82.41552, 79.1805, 78.35847, 78.20818,
  55.77341, 53.28761, 53.70036, 56.36147, 59.49675, 62.47518, 65.53045, 
    68.57973, 72.55824, 76.6787, 80.41323, 83.29762, 85.08586, 86.05365, 
    85.74228, 83.90302, 80.16343, 76.12582, 72.7907, 70.31123,
  56.83235, 61.31199, 66.63993, 70.25359, 71.86951, 72.9725, 72.60254, 
    70.91098, 69.96646, 70.44041, 72.79869, 76.22404, 78.92303, 80.06778, 
    79.95045, 79.00449, 74.78932, 68.97203, 65.02283, 62.69532,
  68.3633, 71.93901, 73.70711, 74.39041, 73.63334, 68.86617, 63.32656, 
    59.99377, 59.12814, 56.99648, 56.24871, 58.72226, 62.77227, 66.22812, 
    68.13854, 68.2399, 66.92085, 65.41513, 64.57212, 64.45194,
  68.09704, 68.24562, 68.24198, 68.9448, 68.36476, 63.28403, 61.62608, 
    61.65208, 62.17025, 60.0423, 54.90421, 56.82523, 64.69385, 70.39545, 
    71.06477, 70.62612, 70.42631, 70.42206, 70.46626, 70.07364,
  90.27865, 90.46936, 90.96187, 91.3328, 91.81367, 92.22416, 92.56532, 
    92.95425, 91.85168, 92.18073, 92.55077, 93.10929, 93.48644, 93.577, 
    93.82186, 94.12104, 93.31866, 93.16252, 93.2915, 93.39014,
  86.08983, 87.35469, 88.52606, 89.70167, 90.95605, 92.19986, 93.32362, 
    94.55434, 91.65786, 92.6256, 93.43529, 94.43275, 95.3866, 96.17465, 
    96.70849, 96.71648, 94.6088, 94.85646, 95.30914, 95.54397,
  86.70512, 88.1973, 89.59498, 90.8068, 92.01413, 93.31496, 94.68686, 
    95.56428, 90.70692, 91.19692, 92.00114, 92.65517, 93.44144, 95.10209, 
    96.78224, 97.73758, 96.97577, 97.40762, 97.64394, 97.73307,
  89.68115, 91.15698, 92.42143, 93.04539, 94.1965, 94.98151, 95.89515, 
    96.40926, 93.8694, 95.00821, 95.94914, 96.63451, 97.44318, 98.08365, 
    98.37001, 98.81956, 99.41076, 99.58131, 99.54997, 99.19375,
  89.67426, 92.05407, 93.37361, 93.45905, 92.23868, 92.88578, 92.82374, 
    92.37224, 90.83638, 91.01794, 91.11318, 91.2873, 91.57444, 91.8625, 
    93.73058, 95.45873, 98.3066, 98.44868, 99.02164, 99.10619,
  85.64087, 88.19569, 89.57105, 89.64063, 89.47247, 89.45906, 88.78096, 
    88.23565, 83.85477, 83.9209, 84.01184, 84.51329, 85.23825, 86.21136, 
    86.95574, 88.00373, 95.86523, 97.04032, 97.85556, 97.95661,
  95.50658, 93.7512, 93.42052, 92.73711, 91.85071, 91.18044, 89.61992, 
    88.19778, 79.25771, 78.88412, 79.78496, 74.28655, 75.03474, 79.51832, 
    82.06604, 79.51465, 86.8036, 90.05141, 92.08651, 92.67957,
  98.3136, 98.21742, 97.58485, 96.61398, 96.4712, 96.65526, 96.51331, 
    96.29932, 91.52852, 91.88051, 92.13867, 88.71255, 87.55116, 91.05211, 
    94.91029, 91.81839, 93.1065, 92.04589, 88.16429, 89.7748,
  97.84018, 97.79051, 97.3247, 97.22118, 97.43619, 97.73954, 98.2092, 
    98.36369, 96.84027, 96.75832, 97.0124, 96.93803, 96.50016, 96.27498, 
    96.29099, 97.09836, 98.19801, 98.8465, 98.63737, 99.01076,
  98.66042, 98.21406, 97.7163, 97.35273, 97.39574, 97.68083, 97.51015, 
    97.31455, 97.22263, 97.32518, 97.31413, 97.33452, 97.54791, 97.75464, 
    97.81731, 98.07378, 98.49442, 98.47986, 98.3119, 98.5476,
  97.26917, 97.16064, 97.05055, 96.79762, 96.50986, 95.69913, 94.08237, 
    93.96456, 94.70052, 94.92776, 95.482, 95.28693, 95.93817, 96.30487, 
    96.15034, 95.95493, 96.05909, 95.82204, 94.18667, 91.53635,
  90.26936, 89.94406, 90.27695, 91.70534, 92.6635, 87.82993, 78.56992, 
    72.90591, 73.91786, 78.82522, 81.69787, 82.86334, 83.01902, 83.81273, 
    87.59975, 88.89301, 89.1429, 86.3702, 77.32833, 70.95148,
  72.60237, 73.85394, 75.07816, 76.11095, 76.13499, 73.10439, 68.69399, 
    66.91071, 67.16811, 68.30428, 69.22557, 70.05745, 71.08477, 73.1063, 
    75.37894, 76.93853, 77.79271, 77.17831, 75.71008, 73.93888,
  70.20754, 69.93935, 69.9543, 70.26144, 69.47583, 67.73914, 66.14673, 
    65.45709, 65.90311, 66.87197, 67.91827, 69.27573, 71.59644, 74.63225, 
    77.81239, 80.20579, 81.0661, 81.54023, 82.13872, 81.50178,
  71.17089, 67.77758, 65.09386, 64.12596, 62.689, 61.44544, 61.04934, 
    61.71202, 63.50428, 65.81725, 68.86181, 72.03522, 74.69347, 76.72852, 
    78.67188, 80.32835, 81.25827, 81.86569, 82.9491, 83.88985,
  70.31931, 65.44547, 60.23208, 58.29305, 57.99087, 58.72477, 60.35605, 
    62.39582, 65.13776, 68.53798, 72.39408, 75.93134, 78.9258, 81.40452, 
    83.10816, 83.79124, 82.47524, 80.27815, 79.85361, 80.03515,
  64.32565, 60.19445, 58.53889, 60.21262, 62.45768, 64.77971, 66.91109, 
    68.5334, 70.27448, 72.38094, 75.34969, 78.60403, 81.39275, 83.18236, 
    83.87424, 83.23768, 80.1152, 76.34571, 73.69403, 71.91177,
  63.61417, 66.56992, 71.09573, 74.41154, 75.77049, 76.05373, 74.96818, 
    72.38411, 69.91143, 68.61705, 68.90154, 70.41422, 72.51038, 74.1751, 
    75.64233, 75.70516, 72.41206, 67.3428, 64.33493, 63.22603,
  74.11085, 77.56428, 78.50999, 78.24831, 77.11918, 72.3632, 66.63581, 
    62.19699, 60.18514, 57.53812, 56.30597, 57.44145, 59.93357, 61.76641, 
    62.72487, 62.82741, 61.81861, 61.21457, 62.44366, 64.02912,
  74.67986, 74.09025, 72.28008, 71.63828, 69.89389, 63.96356, 61.31358, 
    62.05498, 63.04865, 61.57388, 57.85167, 59.0917, 65.77415, 68.85236, 
    68.07928, 67.32264, 67.94349, 69.2151, 71.08256, 72.47744,
  93.04568, 93.01112, 93.33428, 93.64684, 93.54208, 93.79078, 94.11816, 
    94.11546, 92.94925, 93.20354, 93.56378, 93.66265, 94.09669, 94.40761, 
    94.87766, 95.00706, 94.36287, 94.86922, 95.37246, 95.17931,
  87.91546, 89.11015, 90.44867, 91.74315, 92.95021, 94.03472, 94.81275, 
    95.75552, 91.95675, 93.16119, 93.58644, 94.43528, 94.88416, 95.44623, 
    95.52204, 96.00824, 94.04001, 94.6801, 95.47627, 95.61149,
  90.18157, 91.78329, 93.09367, 94.10188, 94.62593, 95.17771, 96.02431, 
    96.81038, 92.01325, 92.94916, 94.26613, 95.76125, 97.00121, 97.3987, 
    96.77382, 96.48228, 96.41441, 97.60815, 98.25105, 99.10908,
  89.8862, 91.50037, 93.05065, 94.16869, 95.1329, 96.11276, 96.99478, 
    97.95014, 95.91473, 97.0166, 97.43277, 97.09196, 97.12125, 97.36758, 
    97.77469, 98.16002, 98.72227, 99.08759, 99.29511, 99.21101,
  87.16335, 88.06263, 89.86611, 91.96803, 93.60877, 94.75459, 95.62978, 
    96.12592, 95.45751, 95.59431, 95.31447, 94.61774, 94.76456, 95.24442, 
    95.91241, 96.32127, 97.86388, 98.25009, 98.61625, 98.90014,
  82.85779, 84.37225, 86.69868, 88.36132, 88.7085, 88.19811, 86.57402, 
    85.14231, 79.98173, 79.8757, 80.10493, 81.35889, 83.3233, 85.50908, 
    87.59556, 90.09531, 97.12043, 98.08211, 98.3543, 98.10835,
  92.87965, 91.47284, 91.66934, 91.03003, 89.63393, 87.53817, 85.16932, 
    84.18885, 75.41856, 75.22541, 76.75064, 69.27393, 71.31108, 79.56635, 
    83.17157, 80.05514, 88.31726, 91.17468, 93.35088, 94.56273,
  96.38414, 96.6512, 97.19339, 96.70306, 96.26802, 96.03889, 94.99522, 
    93.95915, 90.75082, 91.08, 94.089, 90.40166, 91.09087, 95.1616, 97.56213, 
    89.69109, 96.03835, 93.48373, 92.36916, 92.33178,
  95.28132, 95.7337, 96.4422, 96.47005, 96.92366, 96.81229, 96.14042, 
    95.19345, 93.11897, 93.40282, 94.52025, 95.79739, 96.64805, 97.10467, 
    97.7802, 98.46096, 98.72215, 99.31957, 99.39532, 99.14392,
  96.25123, 96.70261, 96.77776, 97.00169, 97.25183, 97.11291, 96.76917, 
    96.57422, 96.02717, 95.6721, 95.51659, 95.65396, 95.56549, 95.71021, 
    95.94229, 96.66721, 96.68552, 97.25195, 97.47217, 97.5812,
  97.5415, 97.52129, 97.1333, 97.13282, 97.39402, 96.9754, 96.70052, 
    96.00925, 94.87958, 94.08837, 94.13777, 93.32083, 92.71771, 92.95763, 
    93.79967, 94.94731, 95.17611, 95.20467, 93.38761, 89.32734,
  96.76878, 96.73467, 96.27477, 95.80989, 95.75227, 94.75697, 90.84474, 
    85.66555, 82.02585, 82.56551, 84.59137, 86.23276, 87.79633, 90.53224, 
    91.97494, 92.57188, 92.95749, 92.15096, 82.43515, 68.9448,
  84.74886, 84.73219, 85.38712, 86.241, 86.41951, 83.87202, 77.38069, 
    71.76228, 68.25037, 66.34049, 64.589, 63.66439, 63.94081, 65.45847, 
    67.23811, 68.84042, 69.20665, 68.13487, 64.41325, 59.2339,
  77.68382, 77.34696, 77.55634, 77.88785, 77.68731, 76.56992, 74.62009, 
    72.57931, 70.86265, 69.83584, 68.80886, 68.26311, 68.3465, 69.3449, 
    70.45822, 70.89925, 69.63084, 69.00183, 69.49906, 69.54823,
  78.47359, 75.68684, 73.58385, 72.6122, 71.1239, 69.54626, 67.85547, 
    66.85558, 67.31096, 69.09978, 71.45095, 74.03161, 76.05937, 77.06158, 
    77.53661, 78.10122, 77.4885, 77.07322, 77.28033, 77.91222,
  76.34395, 73.01936, 68.52595, 65.81129, 64.91156, 64.94664, 65.12791, 
    66.24604, 68.22504, 71.83076, 76.30969, 80.25866, 82.93634, 84.55123, 
    85.12576, 84.82114, 82.72492, 79.86835, 78.8552, 78.89582,
  69.8306, 66.22531, 63.49096, 63.99471, 65.92504, 67.95088, 69.84761, 
    71.61213, 73.31142, 76.14895, 79.67676, 82.76501, 85.00791, 86.56315, 
    86.89462, 85.96016, 82.33929, 78.02926, 74.6761, 72.54919,
  65.47105, 67.41162, 70.88651, 73.25835, 74.43712, 74.60931, 74.31413, 
    72.77502, 70.8173, 71.05651, 72.77186, 74.92172, 77.17539, 79.11314, 
    80.34573, 80.14992, 75.57568, 69.35758, 65.80669, 65.33796,
  74.27321, 75.96491, 75.58652, 75.39233, 74.73765, 72.17835, 68.31049, 
    64.49399, 62.05601, 58.69873, 57.10399, 57.56573, 59.86617, 62.44339, 
    64.7847, 65.87351, 64.89458, 63.79588, 63.78657, 64.84123,
  74.381, 72.08558, 69.73653, 70.15785, 70.00477, 66.96921, 64.7054, 
    61.74247, 62.85329, 61.28238, 57.27003, 56.47181, 60.8853, 64.53764, 
    65.13959, 65.70812, 67.11807, 68.60696, 70.11653, 71.5705,
  91.15371, 91.64606, 91.92358, 92.42795, 92.69508, 93.13999, 93.55474, 
    94.05317, 92.58059, 93.12912, 93.20304, 93.54602, 93.73812, 94.1358, 
    94.36053, 94.50939, 93.83556, 93.86312, 94.07777, 94.07893,
  85.77802, 87.04877, 88.38704, 89.6304, 90.92393, 92.23146, 93.43456, 
    94.53791, 91.27178, 92.17065, 93.13489, 93.92613, 94.7787, 95.51057, 
    96.43332, 97.10088, 95.31227, 96.06112, 96.49048, 97.02405,
  84.40434, 86.15034, 88.10328, 90.00174, 91.74222, 93.37492, 94.69178, 
    95.80022, 91.58699, 92.48892, 93.1506, 93.95843, 94.75599, 95.56576, 
    96.23351, 96.613, 94.75645, 95.03063, 95.40468, 95.79101,
  87.77106, 89.65005, 91.85762, 93.65803, 95.2403, 96.39464, 97.16394, 
    97.83688, 95.76151, 96.22354, 96.24271, 96.39536, 96.60401, 96.88469, 
    96.90741, 96.90664, 97.84052, 97.88377, 97.68481, 97.21042,
  86.84937, 90.20615, 92.95303, 94.68727, 95.69639, 96.285, 96.74591, 
    97.08733, 95.76949, 95.54977, 95.78676, 95.95503, 96.39266, 96.74354, 
    97.016, 96.9723, 99.68557, 99.75405, 99.53229, 99.18038,
  85.65401, 88.83691, 91.37572, 92.86643, 93.63965, 93.85671, 93.52273, 
    93.26603, 88.83273, 88.60059, 88.51091, 88.91911, 89.65063, 90.44458, 
    91.19499, 91.91723, 97.68549, 97.93031, 97.74449, 96.86849,
  93.32104, 91.98441, 92.12479, 91.78726, 92.45681, 92.18958, 91.86021, 
    91.3591, 83.01519, 83.94754, 83.42046, 79.80679, 80.98781, 84.84328, 
    86.3844, 84.96145, 91.22262, 93.00529, 94.2037, 94.55507,
  95.80008, 95.80746, 95.80212, 95.00311, 95.69746, 95.73315, 95.38146, 
    95.21385, 90.37829, 90.29966, 87.39861, 86.20663, 86.29668, 90.37193, 
    93.50173, 84.70405, 92.57561, 92.82619, 91.57355, 92.52868,
  95.59316, 95.63663, 95.59396, 94.67964, 94.27215, 93.84779, 92.84105, 
    92.34722, 90.92516, 91.59765, 91.66474, 91.58811, 91.60677, 91.45694, 
    91.29329, 92.1767, 93.51922, 95.03122, 94.73696, 94.86124,
  96.37835, 96.31588, 96.41499, 96.14897, 95.41566, 94.63109, 93.58985, 
    92.81449, 91.97757, 91.74273, 92.05984, 92.80077, 93.37633, 93.78384, 
    94.33792, 94.54093, 94.79732, 94.77396, 94.61591, 95.01935,
  96.29398, 96.32382, 96.40867, 96.16432, 95.11314, 94.22218, 93.84365, 
    93.68374, 93.00372, 93.40615, 93.3159, 93.16382, 93.30446, 93.6564, 
    94.12247, 94.5186, 94.51991, 94.29578, 94.09801, 94.02351,
  94.31135, 94.27851, 94.06306, 93.13307, 92.28603, 92.05264, 90.23618, 
    87.62183, 86.96881, 88.44827, 88.65465, 88.57573, 88.23403, 88.89684, 
    90.13629, 91.41354, 92.31714, 92.47446, 91.53053, 88.27341,
  85.0923, 83.59087, 82.32201, 80.64777, 79.17335, 77.14263, 73.28564, 
    70.76534, 70.91208, 72.26115, 73.42686, 74.86678, 76.8924, 79.19158, 
    81.38071, 83.43264, 84.64964, 84.71628, 83.17657, 79.0485,
  73.04491, 71.99938, 71.09983, 70.32201, 69.34708, 68.30872, 67.51674, 
    67.63772, 68.23384, 69.62919, 70.9549, 72.98766, 75.83382, 79.09029, 
    81.855, 83.42939, 83.2842, 82.94468, 82.94131, 82.41446,
  73.38241, 70.14858, 67.63133, 66.21286, 64.74073, 63.68108, 63.13287, 
    63.28455, 64.46104, 66.69846, 69.66656, 73.54329, 77.80111, 81.30379, 
    83.46463, 84.28622, 83.96149, 83.40331, 83.77828, 84.6938,
  72.96913, 68.82806, 64.17751, 61.52683, 60.66856, 60.9693, 61.57088, 
    62.78014, 65.63023, 69.3909, 73.55317, 77.67473, 81.16293, 83.97594, 
    85.47735, 85.94878, 85.16603, 83.42224, 82.87695, 82.53791,
  66.43298, 62.33318, 59.67908, 60.63464, 62.82475, 65.04382, 66.96563, 
    68.60876, 70.52805, 72.79861, 76.12594, 79.22063, 81.67229, 83.60358, 
    84.78307, 85.16417, 83.15094, 79.84762, 77.13334, 74.70882,
  63.31979, 64.93928, 69.07435, 72.23227, 73.7208, 74.0975, 73.87026, 
    71.73896, 68.83328, 68.50027, 70.42153, 72.60784, 74.50435, 75.7682, 
    76.57062, 76.68405, 72.97583, 67.94102, 64.92516, 64.55787,
  72.07996, 74.99599, 76.62151, 76.48338, 75.56196, 72.41358, 67.90956, 
    62.75484, 59.04048, 56.81846, 56.3224, 56.8675, 58.03379, 59.31029, 
    60.72761, 61.61808, 60.88291, 60.74584, 62.38142, 64.82382,
  73.26157, 72.64816, 71.84402, 71.78101, 69.9379, 66.24659, 64.30676, 
    62.27598, 63.21777, 62.16458, 59.77563, 57.82189, 61.21847, 63.53283, 
    64.0239, 64.89086, 66.21326, 67.89471, 69.70627, 70.75082,
  90.42122, 90.80277, 91.25312, 91.64415, 92.0071, 92.27158, 92.61368, 
    93.0102, 91.52238, 91.62126, 92.07262, 92.46264, 92.66057, 93.05011, 
    93.36557, 93.19834, 92.43936, 92.60781, 92.85104, 92.9407,
  84.5911, 85.31496, 86.1413, 86.97018, 87.80996, 88.6683, 89.50067, 
    90.37122, 87.02844, 87.99988, 88.98993, 89.98455, 90.96424, 91.98736, 
    92.8723, 93.65512, 91.7242, 92.38094, 92.95825, 93.40704,
  82.75574, 84.23089, 85.76087, 87.13051, 88.38058, 89.63579, 90.84464, 
    91.97983, 87.79185, 89.0823, 90.14006, 91.11827, 92.13338, 93.20409, 
    94.59367, 95.39491, 93.43497, 93.94788, 94.08938, 94.92157,
  83.9454, 86.04388, 88.02225, 89.68379, 90.97329, 92.14191, 93.29279, 
    94.31348, 91.88355, 92.89734, 93.72415, 94.46863, 94.91987, 95.43314, 
    95.69993, 95.79507, 96.41911, 96.14629, 95.97573, 95.8828,
  83.04197, 85.62231, 87.7744, 89.31923, 90.85653, 91.74253, 92.23038, 
    92.91098, 91.60323, 92.34658, 93.09651, 93.57317, 93.97926, 94.37844, 
    94.59666, 94.49812, 97.84132, 97.34921, 96.87173, 96.04736,
  83.84949, 86.51296, 88.35062, 90.2588, 91.32429, 91.52393, 91.51956, 
    91.14906, 86.39048, 86.46471, 86.9073, 87.45026, 88.08546, 89.05531, 
    90.0625, 91.07013, 97.05874, 96.75054, 96.26074, 95.828,
  91.52124, 90.54931, 90.22392, 91.50164, 92.12584, 91.50919, 90.88728, 
    90.61153, 82.85748, 83.86365, 83.93969, 81.37093, 82.50116, 87.24639, 
    88.35151, 86.5319, 92.58073, 94.03619, 94.85804, 94.86945,
  93.85844, 93.90245, 93.83595, 93.87542, 94.18085, 93.79465, 93.26324, 
    92.97941, 88.19899, 88.70315, 86.84979, 86.19001, 87.1401, 91.66802, 
    92.84608, 87.67258, 92.44729, 93.61783, 92.04987, 93.02734,
  94.93122, 94.94533, 94.67984, 94.45795, 94.09769, 93.71172, 93.34532, 
    93.03474, 91.30673, 91.76191, 91.96509, 92.22393, 92.02311, 91.99171, 
    91.93087, 92.69193, 93.03432, 94.986, 93.74834, 93.43693,
  95.50491, 95.17035, 94.86053, 94.7202, 94.64052, 94.2048, 93.71978, 
    93.29131, 93.14043, 93.31482, 93.55454, 93.65807, 93.80347, 93.39631, 
    93.38364, 93.77319, 94.31275, 94.58147, 94.57697, 94.93678,
  95.88468, 95.92992, 95.71816, 95.51121, 95.33961, 95.20732, 95.23055, 
    94.87098, 94.47318, 93.8367, 93.85621, 93.55245, 93.19547, 93.10887, 
    92.96638, 93.16071, 93.32763, 93.38878, 93.54241, 93.91999,
  94.61549, 94.94106, 95.27882, 95.59342, 95.65878, 95.43943, 94.59076, 
    93.6228, 92.8604, 92.42921, 92.10188, 91.53067, 91.06626, 90.64751, 
    90.74429, 90.67, 90.14998, 90.00076, 89.41419, 88.33431,
  91.19661, 91.27988, 91.31909, 91.39619, 91.05535, 89.78207, 86.92182, 
    84.16907, 82.98909, 83.03976, 83.22502, 83.32658, 83.65804, 84.5928, 
    85.87805, 86.8039, 86.50294, 85.88312, 84.09966, 79.78368,
  85.09951, 84.93914, 85.01035, 85.00024, 84.42791, 83.13707, 81.64735, 
    80.73404, 80.70117, 81.42203, 82.02776, 82.92055, 84.35056, 86.2497, 
    88.14723, 89.19019, 87.7689, 86.33771, 85.50678, 84.62518,
  84.97021, 82.53236, 80.68978, 79.70538, 78.34628, 77.1303, 76.26752, 
    76.03555, 76.81287, 78.71999, 80.72459, 82.73605, 84.93163, 86.61477, 
    87.71955, 88.07137, 86.92056, 85.96445, 86.03296, 87.07906,
  82.94598, 79.9345, 75.82194, 74.09995, 74.32117, 75.04804, 75.02963, 
    75.07128, 76.75874, 79.64248, 82.26644, 84.16467, 85.56067, 86.55998, 
    86.66525, 86.55143, 85.80209, 84.86922, 84.84178, 84.68322,
  79.00369, 76.73227, 74.88137, 75.78338, 77.23271, 77.54524, 77.37255, 
    77.67656, 78.74746, 80.30835, 81.67067, 82.81736, 83.77968, 84.42886, 
    84.13789, 84.03044, 82.77343, 80.76899, 78.72489, 76.64574,
  77.0951, 78.49044, 81.31978, 82.89568, 82.71445, 81.47357, 79.45661, 
    76.52807, 74.18031, 74.06038, 74.83857, 76.12494, 77.57824, 78.30867, 
    78.52434, 78.48399, 75.94555, 72.08482, 69.29042, 67.86743,
  80.27109, 82.10825, 81.79823, 80.15726, 79.37558, 77.75469, 73.30666, 
    68.30809, 66.00372, 64.09939, 63.2723, 63.86584, 66.19508, 67.91019, 
    69.45724, 69.5265, 67.47792, 65.84248, 65.78419, 66.64419,
  76.85674, 75.92261, 74.74534, 74.4455, 75.00552, 73.36916, 70.0812, 
    65.2047, 67.09163, 66.51481, 64.61439, 62.50356, 66.61111, 69.46748, 
    68.3384, 67.79736, 67.80563, 68.9177, 70.8996, 72.38713,
  92.79357, 93.07484, 93.258, 92.90774, 93.06613, 93.50137, 93.68522, 
    93.76571, 92.38165, 92.57596, 92.62645, 92.90495, 92.92089, 93.00901, 
    93.29243, 93.53072, 92.5662, 92.76414, 92.67139, 92.81436,
  85.21513, 85.33395, 85.32613, 85.33727, 85.61659, 86.01477, 86.71255, 
    87.28749, 83.67496, 84.37646, 85.20777, 85.85134, 86.23774, 86.7051, 
    87.4756, 88.09651, 86.09753, 86.64458, 87.22385, 87.58643,
  81.23885, 81.1832, 81.05779, 81.13023, 81.67665, 82.0275, 82.50327, 
    83.34995, 79.37698, 80.30883, 81.4035, 82.87122, 84.05641, 85.29722, 
    86.85031, 87.83092, 85.76967, 86.37657, 86.8361, 87.84177,
  81.88297, 82.91073, 83.63583, 83.94405, 83.86859, 84.00191, 84.7067, 
    85.57265, 83.25921, 84.46357, 85.68095, 86.69373, 87.51066, 88.39986, 
    88.82588, 88.86732, 89.77082, 89.53252, 89.20638, 88.98952,
  82.03133, 83.68234, 84.99849, 86.26138, 87.0225, 87.79839, 88.78643, 
    89.75584, 88.56397, 88.90893, 89.54542, 89.97912, 90.13933, 90.2427, 
    90.21241, 89.7132, 94.17902, 93.45422, 92.92005, 92.07182,
  81.69108, 84.03267, 85.59128, 86.65467, 87.39933, 88.19631, 88.50083, 
    89.07713, 85.13365, 85.75121, 86.33511, 86.82621, 87.79581, 88.16807, 
    89.50861, 90.62656, 97.24666, 97.61192, 97.61391, 97.31044,
  87.16315, 84.76291, 84.26799, 84.57947, 84.82309, 84.99268, 85.37115, 
    85.27183, 77.71121, 77.54987, 75.70411, 77.75653, 79.40429, 83.35139, 
    85.89902, 87.48838, 94.54649, 96.32927, 97.39835, 97.67136,
  90.63519, 90.06023, 90.44818, 91.05961, 91.35709, 91.21436, 90.87664, 
    90.46308, 84.03091, 81.76242, 76.41688, 81.71923, 83.56461, 89.33959, 
    89.58858, 81.47697, 83.73679, 92.91259, 92.47585, 94.23307,
  92.54026, 92.07899, 91.62393, 91.24239, 91.19329, 91.40179, 91.35425, 
    90.70581, 88.50974, 88.19982, 87.89048, 87.93823, 88.41982, 89.1162, 
    90.48424, 92.38495, 92.80774, 92.83627, 92.70408, 94.788,
  93.82963, 93.83222, 93.73023, 93.42859, 93.37144, 93.45832, 93.58628, 
    93.78898, 93.83195, 93.52685, 92.715, 91.70871, 91.00614, 90.3836, 
    90.41336, 91.15279, 92.37167, 94.12625, 95.19012, 95.19505,
  93.31054, 93.22653, 93.08261, 92.50187, 91.56213, 91.18214, 91.35011, 
    91.54338, 91.89615, 91.85915, 91.53765, 91.41559, 91.73129, 91.25396, 
    89.4569, 87.47451, 87.12298, 88.5043, 90.01418, 90.93999,
  90.59514, 89.87527, 89.09971, 88.32581, 87.9101, 87.66795, 86.67981, 
    86.16586, 86.8413, 87.66302, 88.44717, 88.76659, 89.0968, 89.28384, 
    88.93222, 87.23588, 86.06339, 86.8313, 87.73507, 87.38585,
  87.07783, 86.85971, 86.7321, 87.02675, 87.35711, 86.79627, 84.29964, 
    81.80209, 80.93963, 81.4426, 81.98756, 82.5825, 83.35999, 84.78716, 
    87.27287, 89.0683, 89.85674, 90.0724, 89.60655, 87.52735,
  85.52457, 84.69917, 83.91556, 83.13712, 82.31325, 81.07169, 79.62166, 
    78.53167, 78.19164, 78.79608, 79.30255, 80.18124, 81.9496, 84.47488, 
    87.5513, 89.91558, 89.78355, 89.28474, 89.56649, 89.463,
  85.83184, 82.93745, 80.35564, 78.92995, 77.62364, 76.82146, 76.55147, 
    76.18568, 76.35037, 77.74653, 79.72871, 81.89265, 84.0993, 85.86676, 
    86.94033, 87.62048, 87.52982, 87.40543, 88.27011, 89.67987,
  82.82246, 80.08652, 77.1691, 76.5509, 77.30361, 78.12787, 77.90356, 
    77.20192, 77.61442, 79.32881, 81.27954, 83.16544, 84.82245, 85.7979, 
    85.9595, 86.2633, 85.95004, 85.43222, 85.98695, 86.18394,
  79.26363, 77.79434, 76.91321, 77.08455, 77.56719, 77.51747, 77.27467, 
    77.25864, 77.49199, 78.18127, 79.15577, 80.32068, 81.4973, 82.44884, 
    83.11741, 83.57356, 82.81762, 81.02629, 79.57153, 79.03866,
  77.84182, 77.34377, 77.46963, 77.13276, 76.62661, 75.95195, 74.91512, 
    72.2857, 69.92699, 69.93441, 70.93331, 72.66975, 74.78707, 76.88239, 
    78.37072, 78.65865, 76.265, 72.71896, 70.88905, 71.50323,
  77.23927, 77.22047, 76.09721, 73.67488, 71.90163, 70.18883, 66.65112, 
    62.32252, 60.39998, 59.78165, 59.83257, 61.0974, 64.39635, 67.6267, 
    69.53103, 69.62187, 68.14825, 67.15332, 68.39189, 70.3014,
  71.9408, 70.27241, 68.58089, 68.74608, 69.79994, 68.76212, 66.15673, 
    61.18927, 62.05839, 62.80636, 63.15414, 62.75204, 65.81199, 69.15247, 
    69.34508, 68.85955, 68.76572, 69.55061, 71.04905, 72.7192,
  92.70583, 92.72906, 92.85115, 93.20866, 93.1391, 93.19375, 93.39628, 
    93.45143, 91.89115, 91.88048, 91.9959, 92.25312, 92.37613, 92.70486, 
    92.79517, 92.81175, 91.88331, 91.99728, 92.20138, 92.44347,
  88.88898, 89.39807, 90.07902, 90.58533, 91.13081, 91.58888, 92.17429, 
    92.76442, 88.96059, 89.44338, 89.94867, 90.45148, 90.97633, 91.51872, 
    92.14496, 92.55653, 90.64331, 91.2428, 91.73222, 92.2587,
  86.30775, 87.08681, 88.38597, 89.5455, 90.64201, 91.58228, 92.7086, 
    93.55463, 89.14814, 90.29137, 90.57678, 90.69044, 91.30821, 91.96011, 
    92.49937, 93.14861, 91.17982, 91.82088, 92.52246, 93.10146,
  85.08212, 86.46973, 87.81398, 88.96862, 90.15485, 91.44592, 92.50375, 
    92.8257, 90.06084, 90.72335, 91.40009, 92.02137, 92.18114, 92.12052, 
    91.66982, 91.15359, 91.3267, 91.06947, 90.98826, 91.25841,
  83.76549, 86.11485, 88.07697, 89.32519, 90.40578, 91.4626, 92.08022, 
    92.39867, 91.15236, 91.60691, 91.75648, 92.10937, 92.07664, 92.23095, 
    92.34636, 92.05728, 96.27563, 95.90228, 95.16777, 94.54259,
  82.27042, 85.11264, 87.29578, 89.04214, 90.43251, 90.76258, 90.99094, 
    91.10733, 86.55244, 86.70856, 87.15236, 88.02512, 89.26795, 90.32475, 
    91.3345, 92.25778, 98.45837, 98.63029, 98.41161, 97.91319,
  87.10021, 84.91785, 84.93576, 85.98331, 86.50809, 86.60345, 86.35571, 
    86.16853, 78.21584, 77.64048, 76.59316, 78.53944, 80.03388, 84.50956, 
    87.7206, 88.48814, 95.45423, 97.15754, 97.75097, 97.82298,
  92.23146, 92.16577, 91.65044, 90.98891, 89.91062, 88.04819, 86.07581, 
    84.25999, 75.89533, 74.47836, 73.7806, 81.18514, 84.0398, 87.48485, 
    77.60973, 75.63035, 78.57562, 94.29065, 94.47697, 96.02266,
  91.2193, 90.40212, 89.72599, 89.59433, 89.33008, 88.58694, 87.39391, 
    86.49968, 83.47099, 83.36198, 83.80383, 84.4919, 85.81435, 87.24565, 
    89.03747, 90.99241, 92.10198, 91.5565, 94.24495, 96.69157,
  90.20242, 89.68059, 89.07819, 89.29986, 89.83372, 90.15658, 89.95894, 
    89.54716, 88.54225, 86.99711, 85.70562, 84.87009, 85.12598, 86.3359, 
    87.90459, 89.34742, 91.47678, 93.48187, 94.89923, 95.02965,
  90.01044, 89.72692, 88.88268, 87.87499, 87.8812, 88.98762, 89.74633, 
    89.68375, 89.79485, 89.35155, 89.0832, 88.92773, 89.23895, 89.2075, 
    88.76626, 88.47148, 89.24776, 89.78516, 90.39549, 90.84927,
  87.72855, 87.37532, 87.44053, 88.1557, 88.67684, 88.82921, 88.39054, 
    88.52185, 89.81778, 90.81558, 91.36176, 91.23718, 90.88681, 90.74982, 
    90.83346, 90.50526, 91.12881, 92.22269, 92.62827, 91.73218,
  89.45244, 89.68774, 89.69378, 89.86064, 89.93679, 89.50417, 87.43844, 
    85.07836, 84.80399, 85.75333, 86.5615, 87.13503, 87.62117, 88.42193, 
    90.0587, 91.7009, 92.87794, 93.02802, 92.88017, 91.33083,
  85.62477, 84.54143, 83.86476, 83.39732, 82.39466, 80.5948, 78.97363, 
    78.43805, 79.59749, 81.47624, 83.08479, 84.82877, 86.63058, 88.63487, 
    90.95786, 92.80032, 93.1731, 92.86739, 92.89964, 92.64547,
  83.07702, 79.38857, 76.75405, 75.47082, 74.00473, 73.18587, 74.15295, 
    76.14993, 78.36121, 80.61633, 82.93502, 84.92791, 86.75276, 88.60899, 
    90.23939, 91.01237, 90.83662, 90.24866, 90.87399, 92.14217,
  78.79999, 75.26179, 72.0584, 71.36671, 72.44469, 74.60607, 77.01754, 
    78.60394, 80.22647, 82.53008, 84.38789, 86.06257, 87.99383, 89.10883, 
    89.08923, 88.59463, 87.46447, 86.7413, 87.92924, 89.02193,
  75.07083, 73.7177, 73.17018, 74.64323, 76.74796, 78.11707, 78.73949, 
    79.14472, 80.20088, 81.37176, 82.62881, 84.10074, 85.38519, 86.05461, 
    85.41919, 84.38893, 82.95277, 82.57442, 83.8847, 85.69988,
  76.48369, 77.38974, 78.89089, 79.75227, 79.93725, 79.57553, 78.21516, 
    74.82092, 71.94337, 72.40543, 74.26749, 76.08146, 77.70051, 78.8651, 
    79.23103, 79.48189, 79.25955, 79.722, 81.31671, 82.88535,
  78.26125, 79.5918, 79.59924, 78.15585, 76.34859, 73.75503, 68.33553, 
    62.06169, 59.75646, 61.04766, 62.9026, 65.1813, 68.03948, 71.03863, 
    73.09583, 75.16939, 77.19022, 78.27455, 78.97375, 79.27312,
  72.79693, 72.769, 71.14326, 69.08615, 68.17456, 66.56525, 65.14984, 
    61.41542, 63.41349, 65.61414, 66.13202, 66.66683, 69.58914, 72.8305, 
    74.20149, 75.70572, 77.11153, 77.89201, 77.05132, 75.83907,
  91.26328, 91.60145, 91.84579, 92.10668, 92.33315, 92.56197, 92.83788, 
    93.0387, 91.52206, 91.82107, 92.25675, 92.61135, 93.00777, 93.37113, 
    93.78864, 93.88147, 93.01225, 93.3584, 93.61464, 93.84084,
  86.96758, 87.72955, 88.51013, 89.22598, 89.94435, 90.89918, 91.7823, 
    92.62855, 89.15443, 89.88326, 90.60005, 91.37135, 92.19009, 93.06493, 
    93.88799, 94.72135, 93.1259, 94.18941, 95.0638, 95.7869,
  86.19858, 87.28941, 88.37048, 89.45456, 90.41154, 91.53922, 92.54251, 
    93.47308, 89.18557, 90.27536, 91.48679, 92.63914, 93.76528, 94.90334, 
    95.87162, 96.77752, 95.03413, 95.54782, 96.12705, 96.78401,
  84.15985, 85.90027, 87.36908, 88.83154, 90.20999, 91.39341, 92.58297, 
    93.67764, 91.41457, 92.82475, 94.21187, 95.03711, 95.72309, 96.47301, 
    97.1405, 97.36044, 98.04243, 97.94881, 97.97694, 97.69524,
  83.26727, 85.76949, 88.02837, 89.59628, 91.23973, 92.66567, 93.59524, 
    94.04115, 92.13865, 92.14246, 92.96667, 94.1391, 95.13073, 95.96074, 
    96.17704, 95.56116, 98.05093, 97.90025, 97.02735, 95.86285,
  82.63007, 85.39271, 87.46679, 89.17599, 90.05942, 90.58632, 90.29137, 
    89.70409, 85.06696, 85.57639, 86.40552, 87.51357, 88.61568, 89.4811, 
    89.83215, 90.34229, 95.88122, 95.76498, 95.63026, 94.85845,
  89.63525, 88.27262, 87.75707, 87.51603, 86.5496, 85.97729, 85.26434, 
    85.65874, 77.94403, 77.74657, 76.60815, 76.27546, 78.76966, 84.18068, 
    87.23457, 83.29222, 89.35817, 91.3289, 92.77951, 93.16802,
  87.01898, 84.50478, 81.8261, 78.38857, 75.34313, 73.46279, 71.56693, 
    70.54421, 63.16817, 62.58971, 63.81389, 72.81225, 75.42923, 81.91115, 
    81.07393, 81.65526, 85.14304, 86.95645, 84.90844, 86.45542,
  82.20783, 81.43171, 80.40063, 79.77774, 78.84322, 77.38066, 75.73199, 
    74.30006, 70.77652, 70.14327, 69.96141, 70.71988, 73.10525, 76.27924, 
    78.95201, 79.72134, 79.18362, 77.55217, 83.825, 88.0265,
  83.35874, 82.85043, 82.32564, 81.69549, 81.18295, 80.72409, 80.22757, 
    79.63129, 79.21888, 78.8965, 78.65776, 79.23164, 80.65341, 82.47045, 
    83.71362, 84.62949, 85.03192, 85.37557, 85.88569, 85.45341,
  87.61831, 87.34454, 87.26519, 86.62285, 85.9207, 85.95735, 85.98182, 
    85.67146, 85.67101, 85.82151, 85.92657, 86.35654, 87.04948, 87.63819, 
    88.4352, 89.33184, 89.95245, 89.87124, 89.57634, 89.13293,
  89.42862, 88.9889, 88.90883, 88.76565, 88.44701, 88.29091, 88.3567, 
    89.00092, 90.23684, 91.64628, 92.5149, 92.47399, 91.88447, 91.54052, 
    91.45772, 91.32801, 91.53257, 91.73484, 91.53756, 90.80643,
  88.39314, 88.44724, 88.45557, 88.50693, 88.57438, 88.37755, 87.63065, 
    87.2239, 87.99855, 89.13181, 90.16599, 91.05843, 91.54522, 91.3706, 
    91.18861, 91.32433, 91.85018, 91.70802, 91.35224, 90.51473,
  83.2769, 82.40056, 81.83305, 81.81855, 81.49155, 80.92557, 80.62244, 
    81.11806, 82.48235, 83.87965, 85.07037, 86.8537, 88.76051, 90.34499, 
    90.79196, 91.12675, 90.47735, 89.87395, 90.03863, 90.12562,
  80.92853, 77.12916, 74.4138, 73.96992, 73.57625, 73.52274, 74.10473, 
    75.61446, 78.04792, 79.94073, 81.98353, 84.32447, 86.44666, 87.87834, 
    88.87703, 89.31812, 89.17209, 88.99256, 89.90827, 91.13013,
  79.03706, 74.40031, 70.30905, 69.57484, 70.71891, 72.4129, 74.32835, 
    76.22193, 78.73299, 81.5993, 83.96099, 85.21662, 86.15022, 87.25639, 
    88.1115, 88.55891, 88.53211, 88.13522, 88.46373, 88.32899,
  74.03026, 72.07845, 71.58685, 72.85542, 74.33098, 75.15328, 75.28473, 
    75.3568, 77.07974, 80.18629, 82.33217, 83.25902, 83.62644, 84.20481, 
    84.29943, 84.11935, 83.37732, 81.84886, 80.56062, 79.5461,
  70.18803, 70.75198, 72.18877, 73.77894, 74.60961, 74.23795, 72.48561, 
    69.3821, 68.26803, 69.95414, 72.37833, 74.36286, 76.28081, 77.2764, 
    78.23228, 78.64809, 76.9935, 74.84343, 74.27042, 75.44029,
  68.87252, 68.90988, 69.73932, 70.2487, 69.5257, 67.25816, 62.43254, 
    57.61004, 56.91596, 58.25465, 59.86382, 62.3505, 66.29232, 70.08858, 
    72.89479, 73.5481, 73.39176, 73.29152, 74.23229, 76.01389,
  65.11118, 64.68005, 63.56782, 62.49925, 62.20929, 60.95686, 59.50586, 
    58.32654, 60.70726, 64.12701, 64.41742, 64.39045, 67.84593, 71.88348, 
    73.36845, 73.93579, 74.26461, 74.48526, 75.02161, 75.71884,
  90.23962, 90.66614, 91.13683, 91.55167, 91.97843, 92.29185, 92.60223, 
    92.95606, 91.7357, 92.11314, 92.41152, 92.72932, 93.12556, 93.5832, 
    94.01425, 94.22498, 93.50925, 93.646, 93.8218, 93.88889,
  85.97031, 87.08288, 88.15931, 89.34943, 90.44781, 91.35188, 92.32027, 
    93.4838, 90.52296, 91.69625, 92.63877, 93.44212, 94.10886, 94.745, 
    95.24244, 95.65135, 93.95591, 94.79914, 95.74892, 96.37549,
  88.84231, 90.57793, 91.96147, 93.04163, 93.73937, 94.48566, 95.02813, 
    95.66689, 91.19154, 92.15147, 93.14037, 94.04124, 94.86369, 95.73912, 
    96.2129, 97.32094, 96.41395, 97.2706, 98.04276, 98.62575,
  87.18143, 88.74137, 90.43748, 92.04164, 93.57539, 94.65493, 95.56763, 
    96.47796, 94.85954, 95.95959, 96.58916, 97.16486, 97.59664, 98.30321, 
    98.87308, 99.24057, 99.62033, 99.64252, 99.54958, 99.16011,
  85.89915, 88.09615, 90.34171, 91.72566, 90.80376, 89.14799, 90.06158, 
    91.34245, 91.45683, 92.75586, 93.05767, 93.9079, 94.88681, 95.86551, 
    96.88954, 97.84422, 99.75259, 99.86357, 99.70674, 99.48833,
  84.6357, 86.1774, 87.03925, 87.75484, 88.13876, 87.71141, 87.29229, 
    86.9258, 82.02043, 81.81429, 82.58743, 84.19396, 85.80888, 87.47978, 
    89.44649, 91.28621, 97.58615, 97.98792, 98.10963, 96.97196,
  92.10596, 90.02838, 89.48897, 90.01364, 89.55316, 89.97391, 90.3751, 
    90.38938, 82.84773, 82.92379, 83.86781, 76.0922, 78.08957, 85.36262, 
    89.40292, 86.13428, 92.95442, 95.17835, 96.1496, 96.15385,
  82.24651, 79.42647, 75.98604, 72.9222, 72.30219, 75.24151, 77.51017, 
    79.18082, 72.83717, 73.99718, 78.44617, 80.26686, 83.46902, 90.60535, 
    93.02876, 94.23264, 94.97993, 93.45391, 88.5794, 88.96692,
  75.96914, 73.6442, 70.91547, 67.92103, 65.13828, 62.86378, 61.23645, 
    60.4471, 58.61827, 58.96691, 59.60195, 60.72873, 64.49291, 69.72006, 
    74.15373, 78.65357, 82.69803, 88.10948, 91.91247, 93.8428,
  81.41633, 81.4401, 81.18076, 79.77778, 77.60808, 75.84695, 74.1852, 
    73.16546, 72.32249, 71.08588, 69.98938, 68.935, 68.32941, 68.10512, 
    67.90612, 68.10161, 68.43636, 70.17178, 72.85571, 75.38261,
  84.09614, 84.52358, 84.77297, 84.02576, 83.11336, 82.43485, 81.73085, 
    81.12797, 80.67327, 79.41838, 77.84908, 76.54546, 75.54516, 75.48005, 
    75.91611, 76.2104, 76.03671, 75.86801, 75.83059, 76.53789,
  84.44726, 84.46062, 84.47896, 84.32672, 83.77056, 82.69624, 81.75839, 
    81.78947, 82.53127, 83.31871, 83.36813, 83.14851, 82.85622, 82.70889, 
    82.63035, 82.52451, 82.59406, 82.1163, 80.76741, 79.14848,
  85.60766, 85.88548, 85.97907, 86.32378, 85.92754, 83.94962, 81.33546, 
    79.66937, 79.92027, 81.76302, 83.11983, 84.14332, 84.96384, 85.42297, 
    85.47267, 85.91467, 86.89213, 87.01991, 85.833, 83.69174,
  81.86817, 81.26277, 81.23256, 81.98635, 81.44608, 79.76859, 78.14055, 
    77.42393, 78.00093, 79.6868, 81.04628, 82.33131, 83.9465, 85.28055, 
    86.11794, 86.86886, 87.18909, 87.08901, 86.87417, 86.18098,
  79.39719, 76.4248, 74.52316, 74.58923, 74.42252, 74.8157, 75.66396, 
    76.89838, 78.24976, 79.88326, 81.55133, 83.21962, 83.99817, 84.06985, 
    84.29522, 84.46224, 83.78383, 82.86688, 83.50984, 85.18552,
  76.00365, 72.94691, 70.08109, 70.23551, 71.77341, 74.22472, 76.52665, 
    78.79829, 80.59871, 81.99361, 82.88532, 83.13961, 82.99202, 82.64651, 
    81.99788, 81.14034, 79.68523, 78.86149, 80.5683, 82.43269,
  71.12182, 70.66351, 71.24512, 72.84848, 74.29401, 75.84637, 77.09703, 
    78.3065, 79.32152, 80.55104, 80.85483, 80.42433, 79.98423, 79.53735, 
    78.66014, 77.20761, 76.05656, 76.18498, 77.27266, 78.70747,
  70.4132, 72.34613, 74.7604, 75.60398, 75.48565, 75.32002, 74.59913, 
    72.40793, 70.34695, 70.00286, 71.03508, 72.41351, 73.54927, 73.8993, 
    73.6927, 73.10992, 72.50108, 72.70144, 74.75037, 76.86505,
  71.50208, 72.74286, 74.15471, 74.06213, 73.43108, 72.06181, 67.65402, 
    62.94106, 60.04227, 58.77795, 59.04659, 60.71129, 63.6751, 66.05376, 
    68.04432, 69.58569, 70.97337, 72.92159, 75.44499, 77.27753,
  67.43958, 68.19278, 68.77596, 68.82707, 68.78732, 68.3681, 67.9866, 
    65.21368, 64.14545, 62.29161, 60.62175, 60.80902, 64.44721, 67.92184, 
    69.98629, 71.80382, 73.80924, 76.31552, 77.73328, 78.16327,
  91.10218, 91.33691, 91.7448, 92.06355, 92.3802, 92.68711, 93.05789, 
    93.52945, 92.26223, 92.77299, 93.25175, 93.77693, 94.45638, 94.88766, 
    95.3068, 95.60217, 95.0359, 95.18687, 95.30954, 95.59646,
  86.04295, 87.48513, 88.99633, 90.52528, 91.98557, 93.45995, 94.43663, 
    96.03044, 93.58707, 94.54686, 95.31512, 96.01735, 96.58019, 96.98485, 
    97.41152, 97.70103, 96.28559, 96.84244, 97.50204, 98.26138,
  86.59929, 88.48552, 90.01505, 91.41861, 92.63615, 93.6359, 94.8268, 
    96.11005, 91.69607, 92.13901, 94.18942, 94.59827, 94.79382, 95.29317, 
    96.05402, 96.33018, 95.88161, 96.42872, 97.72369, 98.49311,
  88.92146, 91.01577, 92.60143, 93.28765, 94.41694, 95.26515, 95.94172, 
    96.63083, 94.28638, 95.55826, 96.69245, 97.48849, 98.09905, 98.47031, 
    99.37157, 99.64746, 99.76804, 99.5511, 99.75886, 99.43724,
  88.27624, 90.76297, 91.62383, 91.40884, 91.73376, 92.22559, 92.75354, 
    93.58809, 93.51062, 94.2999, 95.23765, 96.16912, 96.60524, 96.21706, 
    94.6076, 95.55671, 98.08363, 99.33829, 99.36618, 98.81835,
  84.93897, 87.08147, 88.59217, 89.50323, 90.57263, 91.38445, 91.60539, 
    91.27328, 86.0834, 85.20914, 84.54992, 84.54898, 84.42986, 85.04396, 
    84.16656, 86.36386, 94.06892, 95.98045, 96.67371, 96.87595,
  93.79877, 92.20354, 92.52897, 93.06442, 93.13155, 92.80074, 91.89659, 
    90.83859, 81.44397, 80.92906, 81.7256, 75.32496, 75.31147, 78.53993, 
    83.44725, 79.89444, 86.89452, 89.19134, 90.08098, 89.45848,
  94.40644, 93.60468, 92.01221, 90.1824, 89.28096, 88.936, 87.77091, 
    87.06492, 80.7747, 81.14557, 83.82207, 76.70664, 77.24174, 83.73087, 
    91.27625, 92.01947, 91.36009, 86.95129, 87.02611, 88.00002,
  77.16043, 77.70753, 77.58164, 77.25932, 77.99962, 79.35989, 80.22307, 
    79.76154, 74.05795, 72.12454, 73.44726, 77.13367, 80.77932, 83.03971, 
    82.80767, 84.13297, 88.89143, 94.0657, 95.771, 94.83883,
  79.5489, 81.06141, 82.21872, 82.66743, 82.5457, 82.38547, 82.276, 81.50951, 
    79.8753, 77.74671, 75.76722, 74.34036, 73.32697, 72.20891, 70.76876, 
    71.25594, 71.86124, 75.47375, 79.76184, 83.40431,
  83.61469, 84.93934, 85.67411, 86.08159, 86.05241, 85.88679, 85.84855, 
    85.51792, 85.06121, 84.19904, 83.03889, 81.79874, 80.51408, 79.23853, 
    77.35229, 75.24727, 72.39709, 69.70444, 67.88029, 67.123,
  85.31602, 86.1744, 86.68023, 86.65443, 86.11879, 84.65405, 83.36006, 
    83.40233, 84.43452, 85.16706, 85.02312, 84.58261, 84.03045, 83.51445, 
    82.62949, 81.25288, 79.21162, 76.85336, 73.45178, 70.67882,
  86.46317, 87.17661, 87.20903, 87.05758, 86.57812, 84.75008, 82.32347, 
    80.93388, 81.4472, 82.41821, 83.04288, 83.81099, 84.68514, 85.39324, 
    85.27837, 84.68788, 83.44114, 81.52749, 78.7525, 75.24749,
  83.76808, 82.71766, 81.93383, 81.33125, 79.95594, 78.24799, 77.22868, 
    77.63258, 79.01498, 80.53313, 82.06072, 83.97598, 86.21649, 88.14484, 
    89.13911, 88.60674, 86.39466, 84.91685, 84.02962, 82.08494,
  80.99551, 77.37466, 74.42963, 73.95764, 73.67511, 73.53889, 74.35168, 
    76.35607, 78.93999, 81.29251, 83.5502, 85.98302, 87.94393, 88.94714, 
    88.84982, 88.01795, 86.15815, 84.71523, 84.71815, 84.78029,
  75.96574, 71.92397, 68.57858, 69.90174, 72.88799, 75.70533, 78.71413, 
    82.07619, 84.8683, 86.98844, 87.99342, 88.2129, 88.09957, 87.46091, 
    86.25916, 84.99554, 82.79924, 80.35929, 80.21407, 80.10458,
  69.48017, 68.5275, 70.80183, 76.14439, 80.56021, 83.91552, 86.18864, 
    87.03166, 86.93363, 87.02873, 87.26309, 86.54037, 85.58259, 84.30672, 
    81.80122, 80.02798, 77.05203, 73.91637, 71.81911, 70.43317,
  68.44729, 73.00046, 78.62458, 82.44098, 83.97683, 84.04809, 82.15565, 
    78.81483, 76.47254, 76.23088, 77.07118, 78.04928, 78.03967, 76.52763, 
    74.3813, 72.75715, 69.95869, 67.05577, 65.42706, 65.37254,
  70.54711, 75.67039, 78.48502, 79.70636, 79.51901, 77.56742, 72.97205, 
    68.86353, 67.89292, 66.70293, 65.65451, 65.28458, 66.87194, 68.89133, 
    70.21199, 69.80697, 68.45108, 67.3617, 67.28345, 67.6506,
  70.21245, 72.67511, 72.79373, 72.79866, 72.47855, 71.83384, 71.57173, 
    68.62325, 69.64566, 70.15789, 68.20743, 66.37227, 68.54221, 72.79107, 
    74.15097, 73.62729, 72.39013, 70.96178, 69.92038, 68.68697,
  91.24291, 91.51492, 91.80656, 92.25696, 92.55415, 92.94696, 93.27243, 
    93.61546, 92.08616, 92.47573, 92.80905, 93.16385, 93.51168, 93.8701, 
    94.10838, 94.42045, 93.61897, 93.86024, 93.98495, 93.99657,
  83.19017, 84.75696, 86.37542, 88.27898, 89.99883, 91.6478, 92.84286, 
    94.13712, 91.22202, 92.4841, 93.31296, 94.07009, 95.64669, 96.50546, 
    96.88382, 97.34514, 95.77669, 96.25547, 96.78736, 97.27997,
  82.62064, 84.9577, 87.45427, 89.5442, 91.02836, 92.51169, 93.54543, 
    94.62785, 90.80411, 92.32656, 94.31936, 95.80244, 96.9116, 97.66511, 
    98.02323, 98.05592, 97.46973, 97.93198, 98.22734, 98.5134,
  84.30044, 86.58015, 88.16307, 89.6334, 90.87123, 92.27562, 93.80431, 
    94.95506, 93.91708, 95.35966, 95.86433, 96.98215, 98.33938, 99.19609, 
    99.43986, 98.96798, 98.38985, 98.59414, 98.86684, 98.97144,
  80.60843, 83.25745, 85.71313, 88.00457, 89.34398, 86.7509, 86.8565, 
    86.99136, 87.6215, 89.33054, 91.32175, 93.66722, 95.61736, 97.0096, 
    97.94843, 98.21684, 99.85365, 99.81551, 99.43201, 99.30133,
  79.79315, 80.89395, 82.39717, 83.21438, 83.15479, 83.63288, 84.51611, 
    85.27319, 82.0854, 83.06593, 84.35745, 85.9977, 87.91273, 90.53428, 
    93.1311, 94.63131, 98.91783, 99.41022, 99.67966, 99.1441,
  94.24335, 89.58893, 88.98943, 88.35575, 87.41068, 87.4452, 86.88279, 
    85.6029, 78.0586, 79.19759, 82.77667, 74.90408, 77.57605, 87.00992, 
    90.97014, 87.47959, 94.28318, 96.37685, 96.99891, 96.91367,
  97.7869, 96.44174, 95.16974, 93.53316, 92.90671, 93.19238, 93.25983, 
    93.11655, 89.24776, 91.28969, 94.72459, 90.58023, 92.15145, 96.26788, 
    98.00292, 95.05874, 97.80309, 97.46427, 93.02085, 93.33749,
  98.04691, 97.01868, 96.68943, 96.09394, 94.9405, 95.39569, 96.02383, 
    96.05422, 93.72541, 93.25117, 93.1423, 93.88914, 94.64923, 95.72026, 
    96.0758, 96.6571, 98.2481, 99.16711, 98.97294, 98.74772,
  85.23783, 83.71966, 82.13449, 79.3606, 75.01898, 72.01637, 73.44112, 
    75.69579, 74.8371, 74.17735, 74.85286, 78.3084, 84.50704, 89.38372, 
    91.82255, 92.41219, 93.34556, 94.56844, 95.79861, 96.35236,
  75.09456, 75.94811, 73.95235, 70.29629, 66.01185, 65.18111, 65.59012, 
    66.70393, 67.96695, 69.14999, 70.23162, 71.35372, 72.76005, 74.29909, 
    74.96099, 74.68732, 73.95329, 73.00727, 72.23656, 72.71017,
  69.60658, 69.77961, 70.02598, 70.15862, 70.32481, 69.72, 69.46699, 
    71.00438, 73.93504, 76.41956, 77.52747, 77.93489, 78.15695, 78.41469, 
    78.36654, 77.53332, 76.27955, 74.23557, 70.93802, 68.53922,
  73.53176, 73.96315, 74.08394, 74.72623, 75.70982, 75.77415, 75.07548, 
    74.85136, 76.47321, 78.14274, 79.16055, 79.88667, 80.80963, 82.15269, 
    83.4705, 83.92005, 83.52821, 82.39857, 79.99744, 76.9981,
  73.95226, 73.88821, 74.23331, 75.35759, 75.75262, 75.37286, 74.79714, 
    74.85619, 76.50708, 78.34427, 79.60924, 81.0307, 82.75677, 84.8998, 
    86.65398, 87.11082, 85.7348, 84.51852, 83.89954, 82.52496,
  75.03234, 72.47826, 70.36628, 69.82176, 69.67237, 70.23294, 71.05544, 
    72.31962, 75.18074, 78.12057, 80.78629, 83.68243, 86.52058, 88.43267, 
    89.1117, 88.55165, 86.28055, 84.06924, 83.36463, 83.34492,
  72.74314, 69.61324, 65.88335, 64.90147, 66.505, 69.45499, 72.38078, 
    75.65042, 79.43532, 82.77954, 85.62681, 87.98861, 89.62334, 90.25685, 
    89.28082, 87.59819, 84.75836, 81.93649, 81.40879, 81.28841,
  67.7049, 65.89254, 65.82496, 68.81316, 72.35396, 75.41212, 77.6332, 
    79.4684, 82.02551, 84.45888, 86.80939, 88.38605, 88.56463, 87.84429, 
    85.89172, 83.74192, 80.58745, 77.48254, 75.49717, 74.22018,
  67.63046, 69.72964, 72.94321, 74.60452, 75.28909, 75.19095, 72.96983, 
    69.33365, 67.90176, 69.1404, 72.74494, 76.27174, 78.23178, 78.21909, 
    77.2566, 76.19537, 73.73399, 70.76385, 69.24652, 68.89217,
  69.08975, 70.82407, 70.98613, 69.73814, 69.53085, 67.19176, 62.39187, 
    58.77352, 58.42928, 57.89793, 57.64861, 58.84017, 61.31955, 64.06445, 
    66.2746, 68.01377, 69.24501, 69.86115, 70.80127, 71.65388,
  63.92056, 62.80882, 62.90206, 63.25115, 63.78418, 63.18598, 64.42503, 
    65.55891, 66.00829, 65.85057, 62.29739, 61.14777, 64.61178, 69.04353, 
    71.23333, 72.35414, 73.70236, 74.25558, 74.59425, 74.19263,
  92.04769, 92.49271, 92.62696, 93.24134, 93.57046, 93.64375, 94.1568, 
    94.43604, 92.98032, 93.36012, 93.47273, 93.98, 93.73866, 93.66767, 
    93.96191, 94.00055, 92.86124, 93.01962, 93.35869, 93.2449,
  87.0505, 88.52619, 89.83167, 91.24058, 92.57039, 93.65966, 94.70125, 
    95.32792, 92.22865, 93.44081, 94.263, 95.4112, 95.75277, 96.27509, 
    96.6116, 97.19747, 95.40201, 95.92937, 95.89362, 96.47565,
  83.33563, 84.96598, 86.51751, 88.61928, 90.60663, 92.10301, 93.29102, 
    93.9757, 89.82117, 91.05148, 92.1192, 93.60532, 94.4255, 95.03161, 
    96.15813, 96.95335, 96.70545, 97.7758, 98.48972, 98.50143,
  83.33122, 85.32514, 87.23279, 89.19049, 90.815, 92.01553, 93.12922, 
    93.99279, 92.33205, 92.69753, 92.98908, 93.99078, 94.91756, 95.94033, 
    97.07598, 98.11646, 98.95934, 99.00463, 98.60312, 98.14326,
  79.90779, 82.73194, 84.70699, 86.26005, 87.55669, 87.94726, 88.29334, 
    89.39317, 89.7641, 89.68135, 90.11023, 90.30166, 90.24079, 90.99908, 
    92.2883, 93.80502, 97.19339, 97.7377, 97.86214, 97.912,
  79.15273, 81.29324, 83.01581, 84.49121, 85.31923, 84.49897, 84.17831, 
    84.90837, 81.13043, 81.07038, 81.70722, 82.9921, 84.00454, 85.19116, 
    86.97233, 89.3149, 96.38726, 97.66824, 98.52415, 98.67178,
  93.72746, 89.94603, 88.12878, 87.70174, 86.39043, 85.19697, 84.1895, 
    84.06397, 76.46068, 77.08381, 78.79787, 73.21432, 75.73225, 82.33839, 
    84.95405, 83.41608, 89.83498, 90.87883, 91.95265, 92.22838,
  98.40141, 97.12236, 95.80628, 94.23388, 93.1307, 94.01556, 94.76492, 
    95.81107, 92.16756, 93.56315, 95.92149, 91.58554, 91.69255, 95.23461, 
    95.96117, 88.09775, 93.83067, 95.39704, 89.80833, 90.86625,
  97.51098, 97.30598, 96.74046, 95.65856, 96.3811, 97.0053, 96.85433, 
    96.37172, 93.79633, 93.6463, 95.11237, 96.57742, 97.35103, 96.80966, 
    96.2411, 96.06264, 96.93187, 98.24513, 97.98293, 97.70506,
  95.32316, 94.7637, 94.75218, 94.80445, 94.64569, 93.58469, 91.41145, 
    92.00436, 92.61922, 92.96899, 94.00404, 95.19169, 96.50851, 96.93503, 
    97.05427, 95.79546, 95.44097, 96.52293, 97.3435, 98.56061,
  94.65764, 95.57382, 96.41339, 95.23053, 91.48898, 81.14718, 73.91697, 
    73.5015, 74.98389, 76.31117, 76.89149, 76.99294, 79.17866, 82.09277, 
    82.32072, 81.7177, 82.23177, 79.92741, 73.69515, 73.12149,
  81.13017, 81.10808, 81.39839, 80.32317, 74.12578, 66.12202, 61.66351, 
    62.98935, 66.56539, 69.2123, 70.42229, 70.84436, 71.43883, 71.91003, 
    72.39696, 72.72847, 73.64909, 74.02824, 72.18025, 70.3606,
  69.13066, 69.03074, 68.36698, 67.44797, 66.5521, 65.11891, 63.85455, 
    63.83776, 65.89544, 67.7523, 69.29614, 70.80694, 72.46402, 74.65527, 
    77.0862, 78.62724, 79.74847, 80.05521, 79.23579, 77.71918,
  68.93494, 67.83337, 67.08067, 66.57942, 65.77158, 64.68427, 63.6918, 
    63.26373, 64.24669, 66.11994, 68.04549, 70.32594, 73.2865, 77.40384, 
    81.42778, 83.66179, 83.96056, 83.7875, 83.83755, 83.08416,
  72.00048, 68.19271, 64.86548, 63.01443, 61.32393, 60.07314, 59.77511, 
    60.29033, 62.18331, 65.27204, 68.88824, 72.86168, 76.89766, 80.57303, 
    83.40197, 84.76959, 84.89035, 84.48205, 85.10735, 86.33457,
  72.47428, 67.76675, 61.4062, 58.40565, 57.74007, 58.66154, 60.52586, 
    63.29183, 68.00169, 73.0135, 77.47998, 81.17826, 83.86703, 85.26777, 
    85.73602, 85.65668, 85.00356, 83.92319, 84.45945, 85.29559,
  66.94392, 62.31505, 59.99768, 61.75825, 64.98129, 68.60287, 72.28076, 
    75.61678, 78.95746, 81.87565, 84.31911, 85.85934, 86.73372, 87.02069, 
    86.58606, 85.6213, 83.51057, 81.22473, 79.57344, 78.11187,
  64.25285, 66.21768, 70.01685, 74.00253, 76.32274, 77.3841, 76.01145, 
    72.56757, 70.48271, 70.33141, 72.22417, 75.83593, 78.97495, 79.48288, 
    79.729, 79.4639, 76.3065, 72.39165, 69.9798, 68.64144,
  71.80802, 75.06707, 77.41055, 77.47428, 76.57629, 71.7683, 65.05545, 
    60.88209, 59.64521, 57.70017, 56.66473, 57.64598, 60.62048, 63.63639, 
    65.74047, 66.53188, 66.22398, 65.32883, 65.4156, 66.32365,
  70.58487, 71.98203, 72.41713, 71.94511, 71.10937, 68.26955, 66.57371, 
    66.25936, 65.86909, 62.93818, 57.50283, 57.36659, 62.57587, 67.64169, 
    69.4816, 70.19408, 71.33804, 72.27596, 72.76159, 72.04973,
  93.4754, 93.83453, 94.17703, 94.55048, 94.81233, 95.18404, 95.50739, 
    95.65121, 94.43068, 94.87785, 95.16085, 95.59369, 95.88476, 96.2882, 
    96.39525, 96.78529, 96.13696, 96.27309, 96.44647, 96.65504,
  85.42258, 86.83463, 88.21719, 89.82777, 91.24827, 92.6515, 93.74377, 
    95.01836, 91.78139, 92.87081, 93.65979, 94.5644, 95.06006, 95.72171, 
    96.61175, 97.35105, 95.74934, 96.66016, 97.35493, 98.13977,
  88.59377, 90.49229, 91.99954, 93.27266, 94.23877, 94.90728, 95.55239, 
    96.2522, 91.06496, 92.34336, 93.87013, 94.894, 95.78283, 97.01148, 
    97.59642, 97.75387, 97.48133, 98.15396, 98.45464, 98.79264,
  87.66502, 89.47938, 91.01182, 92.42122, 93.60771, 94.38946, 95.33422, 
    96.41772, 95.24554, 97.14249, 97.85433, 97.94616, 97.74361, 97.68217, 
    98.24388, 98.90162, 99.4444, 99.25026, 98.94553, 98.2287,
  82.24243, 84.78301, 87.25128, 89.56104, 91.37188, 92.15562, 92.53341, 
    93.25629, 93.0771, 93.73563, 94.18842, 94.22968, 94.24527, 94.52701, 
    94.99976, 96.0499, 98.01711, 98.18525, 97.80167, 96.80219,
  81.46418, 83.18897, 84.3297, 85.37285, 86.59341, 87.7641, 87.89799, 
    88.55396, 84.20637, 83.95074, 84.47863, 85.66513, 86.92177, 88.70373, 
    90.21163, 91.46931, 96.67352, 97.08356, 97.39249, 97.46175,
  94.43616, 90.67187, 89.29492, 88.82883, 88.04544, 87.59158, 87.32713, 
    86.97776, 79.93296, 81.04743, 81.91958, 74.53914, 76.94897, 84.42231, 
    86.85342, 85.84666, 92.53053, 94.0947, 94.92901, 95.22658,
  99.03848, 98.5065, 97.75474, 96.85593, 96.8488, 97.20259, 97.06722, 
    97.43761, 94.87665, 95.68083, 95.61303, 93.67432, 94.28915, 96.69456, 
    97.69701, 88.26226, 96.19077, 94.90489, 91.8213, 92.72672,
  97.20039, 97.16828, 97.49591, 97.37792, 97.16404, 96.76015, 97.56513, 
    97.18661, 93.92689, 94.02643, 95.09942, 97.36221, 98.19012, 98.48491, 
    99.00255, 99.18432, 97.38622, 99.71305, 99.01064, 98.59377,
  94.49413, 94.49592, 94.93665, 95.2912, 94.80409, 94.01118, 92.93202, 
    92.18737, 92.41971, 93.3614, 95.09401, 96.48992, 96.81304, 96.36493, 
    95.74524, 95.98064, 96.25899, 97.32879, 97.28713, 97.03169,
  95.09979, 95.34799, 95.35439, 95.02612, 94.87833, 94.09872, 92.30906, 
    91.31197, 90.98102, 91.80174, 92.83763, 93.15422, 93.68304, 93.82955, 
    94.09823, 93.53463, 93.4088, 91.98382, 88.09846, 82.82376,
  92.84781, 93.18594, 93.34753, 93.22681, 92.27502, 87.72198, 78.46327, 
    72.75737, 70.65536, 69.77849, 68.18897, 67.03482, 66.64771, 67.77385, 
    68.84467, 68.26488, 68.99915, 70.31664, 65.154, 62.03901,
  82.25606, 82.30257, 81.81329, 80.58888, 78.98471, 75.08527, 69.65993, 
    65.96957, 64.36827, 63.95269, 63.77375, 63.95161, 65.11271, 66.83494, 
    68.75955, 70.36172, 71.30206, 71.78442, 71.1129, 70.05235,
  80.36685, 79.55965, 78.09605, 76.05904, 73.56917, 70.62545, 68.45354, 
    67.30155, 66.81871, 67.24458, 67.56004, 68.47903, 70.02843, 71.83312, 
    74.00375, 75.49377, 75.46546, 75.45167, 76.28459, 77.10921,
  81.28443, 77.76817, 74.11074, 71.24526, 68.11294, 65.57443, 64.32533, 
    64.47307, 65.24622, 66.30977, 67.97004, 70.52003, 73.132, 75.06065, 
    76.4721, 77.69081, 77.99643, 77.58514, 78.18009, 80.01946,
  79.43561, 74.50008, 67.81782, 63.72218, 62.47141, 62.60964, 63.44919, 
    65.04444, 67.57548, 71.21979, 74.8368, 77.58562, 79.43067, 80.37872, 
    80.2953, 79.4809, 77.68447, 75.72929, 76.25972, 78.06284,
  72.67752, 65.62975, 61.29613, 62.35038, 64.57273, 66.7084, 69.55653, 
    72.80737, 75.8744, 79.13271, 81.61031, 83.31054, 84.08607, 83.49241, 
    81.23109, 79.00861, 75.94167, 72.86498, 71.05573, 70.06973,
  63.43905, 65.0065, 68.92947, 72.09508, 73.59382, 74.21349, 72.64165, 
    69.50308, 67.40457, 67.98201, 70.40112, 73.88706, 76.27477, 75.66225, 
    73.92191, 72.47857, 68.39801, 63.49226, 61.00784, 60.63913,
  68.27464, 72.06697, 73.5787, 73.00114, 71.76627, 67.27808, 61.02493, 
    57.05724, 55.30443, 53.03124, 51.3016, 51.86431, 54.45771, 56.88251, 
    58.57987, 59.1697, 58.69998, 57.97528, 58.88499, 60.87057,
  67.35787, 67.58686, 67.37574, 66.91148, 65.50271, 61.36477, 58.90587, 
    62.73839, 63.6389, 60.86514, 53.33435, 52.01709, 56.49579, 60.8173, 
    62.21513, 62.95658, 63.8308, 64.80383, 66.67517, 68.55505,
  88.71904, 89.0666, 89.46172, 89.9642, 90.48009, 91.05553, 91.5921, 92.146, 
    90.96451, 91.5159, 92.02796, 92.50473, 92.94959, 93.44847, 93.68159, 
    93.93243, 93.23878, 93.44478, 93.65525, 93.82648,
  80.90996, 82.18233, 83.58768, 84.89216, 86.25902, 87.65015, 88.88392, 
    90.08077, 86.91978, 87.88915, 88.70206, 89.38781, 90.13013, 91.14143, 
    91.9832, 92.88799, 91.47026, 92.53476, 93.65778, 94.75821,
  79.53096, 81.68255, 83.85683, 85.9521, 87.77123, 89.35477, 90.91621, 
    92.16835, 87.56769, 89.01246, 91.11476, 92.51405, 93.68093, 94.4707, 
    95.15162, 95.67632, 94.56319, 95.18906, 95.60274, 96.0182,
  80.60196, 83.62003, 86.8607, 89.33092, 91.16885, 92.76718, 94.37144, 
    95.94244, 94.71177, 96.17773, 97.46078, 98.30329, 98.70412, 98.95955, 
    99.11444, 99.24269, 99.60539, 99.53527, 99.21294, 98.83662,
  77.49953, 80.62712, 84.09079, 87.20218, 90.12157, 92.41996, 94.29504, 
    95.66152, 95.97826, 96.48263, 97.01529, 97.10555, 97.6056, 98.08385, 
    98.4528, 98.51333, 99.58444, 99.4992, 99.34837, 98.43314,
  78.06786, 81.09045, 83.87749, 85.99512, 87.24339, 88.28453, 88.7289, 
    89.11014, 85.15305, 85.5034, 86.26189, 87.64484, 89.46574, 91.4913, 
    93.18717, 94.88101, 98.533, 98.64909, 98.92839, 99.16783,
  93.96935, 89.93378, 89.10246, 88.71046, 87.57417, 87.92712, 87.41978, 
    87.65112, 80.48067, 81.17647, 82.11575, 78.11388, 80.39421, 88.02103, 
    89.74142, 87.90002, 93.53676, 94.72692, 95.74206, 96.27238,
  98.77454, 98.54995, 98.18159, 97.66839, 97.25583, 97.69482, 97.57687, 
    98.33128, 95.05209, 94.63374, 95.02879, 94.23782, 94.5017, 96.25961, 
    97.33209, 87.41022, 96.87753, 96.05663, 94.57097, 95.10763,
  96.8065, 97.20007, 96.83575, 96.55521, 96.35834, 97.07992, 97.05681, 
    96.91413, 96.2344, 96.43381, 96.99371, 97.05064, 97.12964, 96.78291, 
    96.63564, 96.90652, 97.25126, 98.73331, 98.54408, 98.5804,
  97.0397, 96.94625, 96.30393, 95.77021, 95.36685, 94.99055, 95.07507, 
    95.83945, 96.52449, 96.79003, 96.99543, 96.81194, 96.71091, 96.75484, 
    96.39484, 96.64758, 96.97128, 97.6953, 98.23337, 97.7421,
  96.53912, 96.99196, 97.0106, 96.60986, 96.35057, 95.86636, 94.8501, 
    93.89926, 93.73795, 94.46787, 95.38654, 95.61505, 95.81711, 96.38572, 
    96.62693, 96.81767, 96.53716, 96.03986, 95.1871, 94.02681,
  93.97415, 93.86769, 93.41658, 93.72238, 94.34746, 93.59896, 91.00797, 
    88.03368, 85.11766, 83.73855, 82.68748, 81.79171, 81.62566, 82.44267, 
    86.40865, 87.91508, 90.14806, 91.29115, 86.8884, 79.85623,
  79.11086, 79.07199, 78.71578, 78.87608, 78.69764, 77.01943, 72.16954, 
    67.1103, 65.451, 65.59113, 65.61574, 65.79921, 67.04462, 69.06351, 
    70.97038, 72.52509, 73.67359, 74.50101, 73.9021, 72.30304,
  72.17233, 71.41061, 70.64042, 69.64365, 67.97083, 66.16202, 64.79034, 
    64.25886, 64.47723, 65.25182, 65.81789, 66.989, 69.12756, 71.88609, 
    74.23413, 75.7254, 75.89551, 75.75999, 76.06795, 76.00043,
  73.72963, 70.78757, 67.79781, 65.84363, 63.84228, 62.28588, 61.62985, 
    61.93087, 63.49532, 65.71874, 67.71655, 70.36108, 73.74044, 76.63931, 
    78.60966, 79.81832, 79.94653, 79.14317, 79.07668, 80.16416,
  72.89226, 69.57762, 64.18522, 60.95368, 60.38438, 60.92553, 62.07866, 
    63.75563, 66.45538, 69.7801, 73.53825, 76.91473, 79.46219, 81.83803, 
    83.35284, 83.4865, 82.16846, 79.56696, 78.78064, 79.45566,
  68.72278, 63.19662, 59.62658, 60.94402, 63.58871, 66.29549, 69.01492, 
    71.58828, 73.99545, 76.83132, 79.67242, 81.70831, 83.04587, 84.17271, 
    84.09528, 82.96336, 80.31348, 77.00234, 74.29365, 71.96101,
  62.07426, 62.81494, 67.04707, 71.10335, 73.2329, 74.3835, 73.78857, 
    71.32201, 69.21264, 69.53218, 71.32914, 74.37684, 76.75418, 78.09402, 
    78.66261, 77.70084, 73.012, 66.96962, 63.10429, 61.22507,
  65.54008, 69.19115, 71.89491, 72.06403, 70.80411, 66.90296, 62.55845, 
    59.61283, 58.2259, 55.99938, 54.52652, 56.20982, 59.17898, 62.04413, 
    64.06214, 64.86462, 63.83706, 62.13748, 61.53144, 61.78527,
  64.77317, 65.71391, 66.19348, 65.85936, 64.38061, 60.748, 59.7023, 
    63.35865, 64.3474, 62.24691, 57.0424, 57.76281, 63.59479, 67.56438, 
    68.30676, 68.69286, 70.21884, 71.51477, 72.21067, 71.95609,
  93.18473, 93.41835, 93.86024, 94.13541, 94.49672, 94.82772, 95.09349, 
    95.48364, 93.97516, 94.40429, 94.73779, 95.16576, 95.47488, 95.74569, 
    96.04818, 96.39091, 95.78316, 96.0141, 96.19501, 96.34348,
  85.6574, 86.94539, 88.311, 89.55965, 90.52288, 91.4749, 92.29123, 93.11443, 
    89.39536, 90.35963, 91.41345, 92.78157, 93.95399, 95.43437, 96.26558, 
    96.83939, 95.71126, 96.74168, 97.50017, 98.02856,
  83.41494, 85.78884, 88.11583, 90.05225, 91.73559, 92.77232, 93.15739, 
    93.25951, 88.94754, 90.73455, 92.79385, 94.46365, 95.78812, 97.04209, 
    97.88791, 98.43873, 97.92664, 98.45991, 98.81491, 99.09287,
  82.91048, 85.40052, 88.43816, 90.80621, 92.26359, 93.31023, 94.43867, 
    95.4129, 94.14036, 95.64626, 97.09624, 98.49961, 99.42129, 99.72377, 
    99.80993, 99.8467, 99.85146, 99.57556, 99.49906, 99.31434,
  80.24473, 82.85383, 85.11411, 86.81808, 89.30047, 91.06853, 92.5408, 
    93.73776, 94.22259, 95.52417, 96.20547, 96.67549, 96.80376, 96.5159, 
    97.28522, 97.83612, 99.35716, 99.37564, 99.37276, 99.43316,
  80.70341, 82.88724, 84.07873, 85.07322, 85.87173, 87.01842, 87.77489, 
    88.34239, 84.54243, 85.25895, 86.15739, 86.88797, 87.63278, 88.47548, 
    89.37711, 90.26675, 96.4862, 97.26379, 97.50478, 97.23915,
  91.27994, 89.55989, 88.7361, 87.98969, 88.06675, 88.41476, 88.30923, 
    87.77768, 79.58772, 79.42683, 79.98766, 75.59544, 76.67979, 81.10452, 
    82.24305, 81.79109, 88.66986, 90.72401, 92.34879, 92.56857,
  96.26445, 96.50409, 96.47786, 96.00199, 96.28954, 97.16733, 97.92907, 
    98.29308, 94.51665, 94.01021, 93.86507, 90.85178, 90.26685, 92.682, 
    94.21763, 84.83716, 91.23316, 88.90665, 88.12995, 89.52145,
  97.03294, 97.24413, 96.78371, 95.7685, 95.23143, 94.89732, 95.07005, 
    94.87008, 92.7261, 94.57312, 95.53061, 96.36082, 96.73213, 97.13712, 
    96.7559, 96.94582, 96.03464, 97.3522, 96.39723, 95.82196,
  96.93353, 97.02463, 96.70819, 95.92078, 94.63573, 93.30637, 93.04354, 
    93.01664, 93.30202, 94.90791, 95.86102, 96.223, 96.23614, 95.81853, 
    96.22758, 97.15449, 97.80287, 98.42627, 98.51614, 98.52453,
  96.71033, 96.60842, 96.40018, 96.16901, 95.65991, 95.05369, 95.5507, 
    95.74954, 95.3326, 95.45067, 95.72993, 96.05586, 95.7483, 95.4163, 
    95.75098, 96.2215, 96.1427, 96.59781, 96.28167, 95.54659,
  96.65619, 96.69091, 96.63638, 96.37489, 95.6019, 94.78458, 94.26707, 
    93.57867, 91.87941, 91.36382, 90.83812, 89.71047, 89.46685, 90.2681, 
    92.32952, 93.0804, 92.90073, 93.43742, 92.02068, 85.64695,
  92.58794, 92.27145, 92.108, 90.948, 88.68244, 85.24072, 81.05573, 78.11077, 
    76.49125, 75.53537, 74.36028, 73.15273, 72.87827, 73.18111, 73.58542, 
    73.68838, 73.31937, 73.52479, 72.70983, 70.03204,
  79.79189, 79.29314, 78.87341, 78.70672, 77.78608, 75.94792, 74.40117, 
    73.54757, 73.34103, 74.10681, 74.75912, 75.62325, 76.83339, 78.05791, 
    78.03818, 77.13219, 75.27022, 74.2932, 74.01398, 74.07172,
  81.15031, 78.96761, 76.55032, 75.42247, 73.78772, 72.06882, 70.83414, 
    70.84695, 71.95853, 74.07137, 76.35632, 78.07997, 79.52341, 80.53172, 
    80.40559, 80.00922, 78.96095, 78.2414, 77.95823, 78.77831,
  81.8195, 79.60789, 74.50011, 71.10043, 69.86823, 70.00775, 70.6433, 
    71.97178, 73.94495, 76.27763, 78.37644, 80.26202, 81.75711, 82.93114, 
    83.45753, 83.44048, 81.74239, 79.30438, 77.9953, 77.69436,
  77.21722, 73.5181, 69.81235, 70.39718, 72.58138, 74.46783, 76.60181, 
    78.78408, 80.21176, 80.95415, 82.20531, 83.50039, 84.34659, 84.66266, 
    84.33043, 83.25063, 79.97825, 75.87863, 71.7436, 68.58717,
  69.75837, 71.57311, 76.44507, 80.70802, 82.80388, 83.8858, 83.86449, 
    81.00132, 77.59939, 76.49303, 77.3371, 78.15049, 79.40022, 79.21213, 
    78.36341, 76.73752, 71.05084, 63.60755, 58.03215, 56.28445,
  77.91764, 81.84052, 84.13726, 84.81001, 83.60319, 79.51188, 73.64592, 
    67.23601, 63.65115, 60.08296, 58.69899, 59.43102, 61.16323, 62.08882, 
    62.22192, 60.8568, 57.21086, 54.73055, 54.58582, 56.51323,
  82.40507, 81.73931, 80.26792, 80.14289, 77.69573, 71.94565, 67.36851, 
    62.10333, 62.39094, 60.10313, 57.66487, 57.62714, 62.56674, 63.88177, 
    62.31284, 61.34711, 61.23783, 62.0337, 63.60153, 65.88108,
  89.33743, 89.6899, 90.14959, 90.61353, 90.99582, 91.40112, 91.80436, 
    92.14952, 90.62619, 90.93166, 91.23126, 91.45008, 91.65788, 91.8343, 
    91.90362, 92.05591, 91.18085, 91.3086, 91.58113, 91.72197,
  83.34271, 84.35603, 85.39888, 86.49144, 87.64915, 88.85686, 90.08018, 
    91.2978, 88.06984, 89.12694, 90.25305, 91.29852, 92.28522, 93.16634, 
    93.8997, 94.49941, 92.58978, 93.2578, 93.78377, 94.30668,
  81.38478, 82.86247, 84.31787, 85.75341, 87.2471, 88.70986, 90.25825, 
    91.60431, 87.52467, 88.9437, 90.48451, 91.93484, 93.13106, 94.11681, 
    95.17325, 95.97296, 94.99854, 95.85117, 96.47988, 96.89296,
  81.1591, 82.79865, 84.58844, 86.69811, 88.80666, 90.76855, 92.52787, 
    94.1153, 92.32034, 93.74942, 95.29098, 96.41039, 96.85693, 97.25404, 
    97.84711, 98.0004, 98.70143, 98.61568, 98.25516, 97.92473,
  78.46672, 80.49895, 82.27342, 83.39826, 84.97202, 86.39605, 87.9554, 
    89.57307, 89.74867, 91.03317, 92.34011, 93.28223, 94.20792, 94.90424, 
    95.46811, 95.73288, 99.24294, 99.18375, 99.04175, 98.25187,
  76.0145, 77.68612, 79.35321, 80.82686, 81.92994, 82.82776, 83.4332, 
    83.94999, 80.3109, 80.76566, 81.4243, 82.37448, 83.62694, 85.11915, 
    86.69302, 88.35394, 95.82899, 96.42381, 96.35052, 95.19209,
  87.69982, 85.33133, 84.97263, 85.0671, 84.83653, 84.53214, 84.92548, 
    84.47581, 76.94516, 78.11326, 79.4466, 74.79231, 76.72341, 83.14639, 
    85.37675, 84.39673, 91.09966, 92.8054, 93.75574, 93.81113,
  92.90674, 93.39281, 94.45874, 94.18504, 94.71486, 94.10635, 95.18098, 
    95.12505, 90.18465, 90.89864, 90.77278, 88.71421, 90.0406, 93.54565, 
    95.69398, 83.21734, 94.64079, 95.69743, 95.23474, 96.06865,
  94.84389, 94.56154, 93.98471, 93.30563, 93.07119, 92.4234, 91.99986, 
    92.04476, 90.90355, 91.54748, 92.05257, 92.57288, 93.05364, 93.19878, 
    93.83727, 94.80613, 95.59969, 96.97606, 96.17978, 96.86403,
  95.3786, 95.188, 94.87141, 94.51458, 94.51762, 94.51206, 94.43328, 94.1458, 
    94.06145, 93.82964, 93.60771, 93.46796, 93.49938, 94.10217, 94.5841, 
    95.05334, 95.74317, 96.33214, 97.02899, 97.14212,
  94.97997, 94.81407, 94.54187, 94.22549, 94.38575, 94.60267, 94.75066, 
    94.90584, 94.96114, 94.9651, 94.65247, 94.24747, 94.50364, 94.84131, 
    94.99262, 95.42284, 95.44685, 95.24462, 95.09952, 94.90986,
  94.40383, 93.76332, 92.90012, 92.70216, 92.47225, 92.42416, 91.47188, 
    90.50835, 90.29465, 90.60612, 90.61454, 90.50554, 90.68126, 91.12893, 
    91.8603, 92.06876, 91.40717, 91.36833, 91.16351, 90.274,
  85.98679, 85.07455, 84.56265, 84.65608, 84.2535, 82.36342, 78.76818, 
    76.45616, 76.58498, 77.48373, 77.93317, 78.45004, 80.01889, 82.39944, 
    84.08618, 84.36626, 83.20786, 81.23363, 79.33215, 77.08048,
  79.27042, 78.59019, 77.86862, 78.11208, 77.50948, 75.82636, 74.39255, 
    73.71155, 73.97707, 74.95485, 76.12056, 77.63366, 79.90121, 82.42058, 
    84.21191, 84.76559, 83.84518, 82.47575, 81.82448, 81.3251,
  81.69385, 79.43264, 76.78022, 74.9017, 72.52785, 70.66381, 69.8297, 
    70.1935, 71.67063, 73.99018, 76.3724, 78.9228, 81.30749, 82.98728, 
    83.44641, 83.49872, 83.08672, 83.04655, 83.60693, 85.02307,
  80.13634, 77.56052, 72.39501, 68.27819, 66.75742, 67.25912, 68.91729, 
    70.85203, 73.45245, 76.17443, 78.69566, 80.76107, 82.49564, 83.69159, 
    83.99081, 84.24255, 84.12298, 83.47017, 83.3401, 84.21685,
  73.63741, 69.6399, 65.54585, 65.38223, 67.45193, 69.95189, 72.51434, 
    74.76379, 76.7049, 78.33539, 79.69836, 80.73174, 81.67593, 82.54086, 
    82.78243, 82.73974, 81.34283, 79.70362, 78.38418, 77.66527,
  67.12714, 67.7604, 71.49389, 74.51753, 75.78526, 76.4871, 76.66041, 
    74.66991, 72.57925, 72.4748, 73.62354, 75.01899, 76.28564, 77.30508, 
    77.56017, 77.04617, 74.60099, 71.41341, 69.29411, 68.673,
  74.37507, 78.41054, 80.92729, 80.60802, 78.63735, 74.81702, 69.94366, 
    65.86303, 63.31497, 60.70046, 60.48775, 61.67748, 64.20331, 66.20415, 
    67.09158, 66.60446, 64.95332, 63.80751, 63.83866, 65.17379,
  77.36516, 78.03805, 77.65268, 76.79948, 75.13847, 70.93074, 67.21999, 
    63.35556, 63.64125, 63.54379, 63.50576, 63.56495, 68.65157, 69.83798, 
    68.06207, 66.54877, 66.01632, 66.45395, 67.67004, 69.34978,
  91.03164, 91.28097, 91.61752, 91.95973, 92.22754, 92.56672, 92.79098, 
    93.0113, 91.5333, 91.80436, 92.14737, 92.36164, 92.66302, 92.44974, 
    92.74084, 93.00687, 92.13474, 92.65121, 92.53175, 92.29919,
  86.45543, 87.15771, 87.89254, 88.64736, 89.36244, 90.24338, 91.06424, 
    91.83907, 88.16501, 88.90138, 89.57915, 90.28169, 90.94241, 91.60615, 
    92.2869, 92.98795, 91.01669, 91.52386, 92.15881, 92.80897,
  86.454, 87.59232, 88.67828, 89.88871, 91.05972, 92.30885, 93.50959, 
    94.58562, 89.97404, 90.70628, 91.38651, 91.98544, 92.62484, 92.88599, 
    93.50397, 94.24358, 92.33147, 92.95686, 93.78066, 94.64265,
  86.38911, 88.026, 89.68391, 91.17489, 92.40681, 93.58733, 94.8343, 
    95.91957, 93.10686, 93.96187, 94.41183, 94.98235, 95.37806, 95.72152, 
    95.91048, 95.9792, 96.79117, 96.71494, 96.67774, 96.77288,
  84.36308, 86.38922, 88.21542, 89.97388, 91.44038, 92.32247, 92.96732, 
    93.26849, 91.83308, 92.17873, 93.05903, 93.99199, 94.67414, 95.2039, 
    95.41373, 95.36415, 98.6088, 98.20151, 97.61953, 96.78014,
  82.83844, 85.85513, 87.95655, 89.50515, 90.74166, 91.523, 91.66437, 
    91.39295, 86.64836, 86.68369, 86.8973, 87.45507, 88.26592, 89.37173, 
    90.56412, 91.45541, 97.28247, 97.33936, 97.09261, 96.2449,
  87.73516, 86.69996, 86.5608, 87.49147, 88.00562, 87.98104, 87.74397, 
    87.37967, 80.20707, 81.04887, 80.55627, 79.37921, 80.86521, 85.09348, 
    85.66039, 85.57058, 91.53709, 93.08141, 94.05972, 94.32873,
  90.23829, 90.73328, 91.21187, 91.69006, 91.73869, 91.54958, 91.84187, 
    92.14884, 86.86732, 86.5873, 82.86548, 83.48249, 83.89099, 87.90614, 
    87.3313, 80.32016, 86.899, 90.82205, 90.70295, 92.09869,
  93.60128, 93.25461, 93.42822, 93.85513, 93.97815, 93.75624, 93.50208, 
    93.6701, 92.00517, 91.71632, 91.42417, 91.04822, 90.99522, 90.33051, 
    90.16823, 90.12318, 89.66879, 90.03291, 88.45037, 90.32394,
  94.48168, 94.42733, 94.51466, 94.63229, 94.93159, 95.05129, 94.80539, 
    94.81108, 95.26125, 95.46204, 95.90756, 95.79111, 95.48862, 95.16948, 
    94.56003, 94.2349, 93.6684, 92.91241, 92.65779, 92.76575,
  93.64377, 93.45482, 93.51498, 94.1236, 94.46765, 94.46847, 94.60721, 
    94.35153, 94.05666, 94.05506, 93.99489, 94.2141, 94.2161, 94.63215, 
    95.01568, 94.83033, 95.02346, 94.79313, 94.30516, 93.59941,
  90.34301, 90.22119, 90.86449, 91.91863, 92.59849, 92.97124, 92.77367, 
    91.68233, 89.90132, 89.36376, 89.22382, 89.98881, 90.57137, 91.22919, 
    91.63299, 91.26761, 91.20918, 91.54472, 90.63564, 88.69952,
  81.18159, 82.18935, 83.20338, 84.39983, 85.04195, 83.34638, 78.58712, 
    75.32941, 75.09383, 76.10467, 76.64239, 77.3367, 78.94695, 82.37279, 
    85.01839, 85.50175, 84.78102, 84.71638, 84.61388, 83.45349,
  77.70988, 75.10642, 73.30026, 72.7862, 71.62514, 69.82963, 68.3576, 
    68.07929, 68.85526, 70.59711, 72.56136, 74.72649, 77.11575, 80.36718, 
    83.81327, 85.05261, 83.85504, 83.40464, 83.88542, 84.64262,
  78.3172, 73.70877, 69.28716, 66.7562, 64.40498, 62.59754, 62.39022, 
    63.85616, 66.2661, 69.61164, 73.31822, 77.32272, 80.53368, 82.88496, 
    84.31273, 85.02184, 84.70762, 84.9175, 86.08461, 88.06949,
  77.0389, 72.65115, 66.49445, 62.22723, 60.63084, 61.17995, 63.31984, 
    66.45231, 69.77917, 73.81361, 77.87593, 81.18223, 84.01479, 85.748, 
    86.07027, 86.29877, 86.11855, 85.55041, 85.27063, 85.31348,
  74.24203, 69.19167, 64.62054, 64.36281, 65.67953, 67.61899, 70.16725, 
    72.64315, 74.94654, 77.21776, 79.67608, 81.67824, 83.30663, 84.5863, 
    84.9636, 85.03011, 83.68312, 81.25957, 78.55561, 76.2393,
  72.16353, 71.67516, 74.39134, 77.47516, 78.77465, 79.5111, 79.03678, 
    75.71975, 71.03969, 69.71835, 71.3148, 74.30459, 77.56703, 79.5259, 
    80.51247, 80.15058, 76.45805, 70.8054, 67.18886, 66.27489,
  75.64956, 78.52003, 81.46165, 82.76732, 81.90303, 79.3966, 74.40202, 
    68.18243, 60.95269, 56.30797, 55.57796, 57.87797, 62.28678, 67.15103, 
    69.96083, 70.45556, 69.00925, 67.28522, 67.27696, 68.75368,
  75.43442, 76.05756, 76.57041, 77.07708, 76.21076, 72.56445, 68.5047, 
    63.25798, 59.40269, 56.30353, 55.99892, 57.904, 65.48466, 71.59864, 
    73.27464, 74.04219, 75.09724, 76.00842, 77.06165, 78.16938,
  92.62572, 92.87477, 93.13387, 93.40256, 93.72988, 94.02205, 94.2672, 
    94.43237, 92.89291, 93.12108, 93.25138, 93.38231, 93.61126, 93.54545, 
    93.78857, 94.00249, 93.20338, 93.30951, 93.36291, 93.55066,
  84.38592, 85.12975, 85.97503, 86.78351, 87.64721, 88.61515, 89.42207, 
    90.22615, 86.97729, 87.85419, 88.86221, 89.85745, 90.69267, 91.31274, 
    91.83704, 92.61418, 90.58128, 90.99089, 91.21751, 91.53719,
  80.55997, 81.6187, 82.90531, 84.15871, 85.33762, 86.75328, 88.14629, 
    89.37418, 85.15607, 86.27068, 87.27205, 88.27684, 89.21216, 90.51756, 
    91.69434, 92.70438, 90.45625, 91.08837, 91.64878, 92.18252,
  79.58333, 81.14864, 82.93066, 84.60998, 86.27402, 87.66496, 88.59937, 
    89.69041, 86.8912, 87.95982, 88.42966, 89.26998, 89.9631, 90.16092, 
    90.69798, 91.03185, 91.8796, 91.72359, 90.89203, 90.46238,
  81.27869, 83.51846, 85.38655, 86.72337, 87.65806, 88.21964, 88.35649, 
    88.54109, 86.73111, 87.16138, 87.69844, 88.06959, 88.14066, 87.94286, 
    88.10636, 87.72036, 92.8227, 92.58912, 91.78926, 90.80302,
  82.23608, 84.88454, 86.80707, 88.0237, 88.70967, 89.06223, 89.02444, 
    88.91233, 84.47909, 84.72712, 85.28368, 86.2836, 87.1228, 87.69151, 
    88.24503, 88.19744, 94.36574, 94.46237, 94.43331, 94.11676,
  87.60294, 85.59511, 85.4134, 86.07663, 86.19493, 85.72894, 85.25964, 
    85.15114, 77.67982, 77.52218, 75.64716, 77.8446, 79.32913, 82.28049, 
    84.04327, 84.40154, 90.50689, 91.86197, 92.76913, 93.4663,
  91.25948, 91.75277, 91.82345, 91.74986, 91.60571, 91.08862, 90.62904, 
    90.34478, 84.60276, 83.04688, 77.28098, 80.77901, 82.08565, 86.81707, 
    87.91332, 82.03088, 84.17574, 90.2375, 88.68492, 90.12281,
  93.27106, 93.40038, 93.40652, 93.32364, 93.35958, 93.48284, 93.53805, 
    93.37952, 91.33153, 91.49542, 91.78304, 91.51381, 91.26011, 91.22191, 
    91.25426, 90.94481, 90.31303, 87.52287, 86.94308, 89.46681,
  93.72826, 93.9826, 93.81049, 93.58672, 93.02816, 92.76867, 92.46161, 
    92.48213, 93.00453, 93.52412, 94.13007, 94.22943, 94.30372, 94.67223, 
    94.80873, 94.80283, 94.34667, 94.07409, 93.48529, 92.82103,
  91.30781, 91.71265, 91.927, 92.08401, 91.6851, 90.99953, 90.85574, 
    91.12344, 91.56889, 91.21522, 90.99624, 91.23692, 92.02602, 93.15876, 
    93.98617, 93.59729, 93.00624, 92.31453, 91.11363, 90.1129,
  87.23492, 87.63606, 88.69857, 89.59157, 90.26398, 89.98401, 89.32961, 
    89.17812, 88.94569, 88.13565, 87.49892, 88.05474, 89.75908, 91.47031, 
    92.44577, 92.91836, 92.56703, 91.40242, 88.94244, 86.523,
  88.76868, 88.55422, 88.89142, 89.53811, 89.35495, 87.57262, 84.34761, 
    81.95408, 81.55356, 81.91135, 82.45205, 84.27527, 86.95754, 89.27744, 
    90.36448, 91.20327, 91.55247, 90.69625, 89.05181, 86.71323,
  87.45101, 85.70428, 84.5345, 84.01614, 82.50531, 79.95651, 77.81738, 
    76.91148, 77.18439, 78.32337, 79.5246, 80.52446, 82.35175, 84.80022, 
    87.08285, 87.94924, 87.25331, 86.35719, 86.33508, 86.12024,
  86.0612, 82.84039, 80.06281, 78.77739, 76.90326, 75.17671, 74.79057, 
    75.60274, 77.14713, 78.77872, 80.18024, 81.82264, 83.30062, 84.14932, 
    85.42023, 86.5309, 86.59457, 86.15807, 86.58962, 88.02082,
  83.50843, 80.45433, 76.25483, 74.06078, 73.27681, 73.67715, 75.55487, 
    77.91324, 80.6321, 82.73536, 84.0448, 85.03394, 85.68456, 86.11607, 
    86.55065, 87.26894, 87.52003, 87.40895, 88.12331, 88.95005,
  78.91055, 75.96642, 72.44361, 72.05608, 73.74168, 75.5808, 77.30567, 
    79.23503, 81.04423, 83.03707, 84.22142, 84.67382, 84.70187, 85.03378, 
    85.60724, 86.52565, 86.50472, 85.86571, 85.18515, 85.2679,
  75.17509, 73.39148, 73.80116, 75.58472, 76.66517, 77.37955, 77.4274, 
    76.02151, 73.99651, 74.2387, 75.89295, 77.90361, 79.63412, 81.00914, 
    82.11852, 82.74923, 81.25233, 78.21503, 76.67453, 77.20649,
  73.12216, 73.72042, 74.04329, 73.72401, 73.09086, 71.62672, 69.03576, 
    65.55053, 61.40323, 58.67473, 58.11934, 60.84002, 66.07968, 70.54962, 
    72.66146, 72.71555, 71.35201, 70.63377, 71.65504, 73.07262,
  69.69509, 68.35408, 67.36819, 67.28154, 67.53863, 65.53922, 62.64829, 
    58.05632, 56.07458, 55.15796, 55.7697, 59.24729, 66.51874, 71.29867, 
    71.54913, 71.03627, 71.03108, 71.94553, 73.828, 74.25826,
  92.92564, 93.14806, 93.42696, 93.68404, 93.91962, 94.07684, 94.26083, 
    94.4565, 93.11724, 93.37776, 93.58154, 93.78804, 94.03655, 94.24667, 
    94.33662, 94.49567, 93.43404, 93.74255, 93.75603, 93.82291,
  86.139, 86.60515, 87.32337, 88.14129, 89.04366, 89.98837, 90.57925, 
    91.41451, 88.21118, 88.78764, 89.54964, 90.36505, 90.75597, 91.51027, 
    92.1199, 92.74394, 90.91013, 91.26971, 91.49422, 92.01154,
  83.20729, 84.18126, 85.18593, 86.23172, 87.20171, 88.21822, 89.15403, 
    90.1628, 86.1129, 87.1681, 88.22795, 89.18254, 90.30568, 91.29362, 
    92.18975, 93.09308, 91.28911, 91.9936, 92.84306, 93.0712,
  83.89709, 85.59076, 86.62768, 87.77552, 88.8494, 89.75357, 90.62057, 
    91.39909, 88.58913, 89.43999, 89.98411, 90.57166, 90.88825, 91.26151, 
    91.84435, 92.06491, 92.9584, 93.63245, 93.98756, 94.28948,
  84.18081, 86.16316, 88.34549, 89.48678, 90.13564, 91.19115, 91.65099, 
    91.94025, 90.42744, 91.07625, 91.36615, 91.68443, 91.92711, 91.9413, 
    92.04135, 92.21871, 96.70943, 96.64523, 96.43306, 96.23057,
  83.72672, 85.95106, 87.52583, 88.81939, 89.97847, 90.47252, 90.95387, 
    91.24022, 86.8391, 87.11195, 87.62807, 88.21334, 88.86031, 89.87125, 
    91.27901, 92.44669, 98.45345, 98.63551, 98.43393, 97.96113,
  88.91055, 86.0547, 85.16903, 85.69044, 85.99608, 86.05182, 85.96393, 
    85.61502, 77.75172, 76.67236, 75.00044, 77.01299, 78.95913, 83.65873, 
    86.48275, 87.67002, 95.04016, 96.82327, 97.8366, 98.07616,
  92.47279, 93.14922, 92.80783, 92.38421, 91.52305, 89.89094, 88.4556, 
    87.36083, 80.82705, 78.83447, 76.53487, 83.34758, 85.00301, 88.47127, 
    83.63088, 80.44799, 85.16066, 92.40426, 92.17253, 93.53748,
  88.15891, 86.9331, 85.48118, 83.69347, 82.77776, 83.15126, 84.06776, 
    84.92242, 83.88541, 85.72476, 87.26251, 88.20538, 89.32011, 89.93955, 
    90.15986, 89.87584, 89.85675, 89.814, 92.57172, 95.34295,
  88.43484, 87.78725, 86.16113, 83.74043, 82.17479, 81.74992, 82.25927, 
    83.08769, 84.29337, 85.42973, 86.76841, 88.07597, 89.19, 89.78298, 
    89.91391, 90.1196, 90.58709, 90.48777, 90.54873, 91.22018,
  87.79279, 87.85771, 86.8604, 85.40718, 84.92367, 85.31801, 86.09495, 
    86.60931, 86.90997, 86.55619, 86.15047, 86.27724, 87.85771, 89.14861, 
    89.75634, 89.48331, 89.48134, 89.28529, 89.21223, 89.27132,
  87.31789, 87.65279, 87.57767, 87.72043, 88.26453, 88.76003, 88.6967, 
    89.155, 89.56026, 89.37699, 88.40101, 87.40329, 87.72031, 88.62234, 
    89.52988, 90.58915, 91.8474, 92.08244, 91.1547, 90.12524,
  88.23763, 88.31981, 88.10595, 88.23789, 88.3023, 87.06553, 84.34332, 
    82.80704, 82.64577, 82.69537, 82.23661, 82.47742, 84.14645, 86.53075, 
    88.69958, 89.84208, 91.07381, 91.81326, 91.85409, 90.95389,
  85.86915, 84.12791, 83.0151, 82.83844, 81.75422, 79.76747, 78.13165, 
    77.22594, 77.28532, 77.99092, 78.37098, 78.90584, 80.65997, 83.36642, 
    86.07629, 87.26132, 87.15216, 87.55098, 88.57515, 89.21084,
  84.7718, 81.06129, 78.54852, 78.45286, 78.0738, 77.28562, 76.63292, 
    76.66708, 77.61476, 79.12304, 80.55389, 82.37267, 84.24222, 85.04122, 
    84.86169, 84.79836, 85.19656, 85.64907, 86.65476, 87.5913,
  82.95587, 80.14877, 77.15878, 76.80717, 77.66035, 78.36048, 78.86679, 
    80.00245, 81.72752, 83.55798, 84.69321, 85.96711, 86.9203, 87.01139, 
    86.19179, 85.47747, 84.86073, 84.35799, 84.35689, 83.54041,
  80.49435, 79.51139, 79.2524, 79.48923, 80.40471, 80.9237, 80.98357, 
    81.4827, 82.26517, 82.86146, 83.74509, 85.03392, 85.98208, 86.2218, 
    85.62314, 85.02358, 83.0284, 81.14239, 79.33386, 76.95956,
  79.53527, 80.2226, 81.18445, 81.5555, 81.46244, 80.7687, 79.69151, 78.2599, 
    77.1479, 77.19711, 78.8017, 81.12883, 82.63799, 83.69958, 83.49717, 
    82.44864, 80.01619, 76.78847, 74.06044, 73.33162,
  76.72205, 76.99213, 76.34472, 75.5202, 75.40344, 74.93951, 73.50534, 
    70.76733, 67.78928, 66.64872, 65.88866, 67.2067, 70.4846, 73.33239, 
    74.2774, 73.19521, 71.50397, 70.85245, 70.6892, 71.13319,
  69.13016, 67.50374, 67.28152, 69.4579, 72.24056, 71.54641, 69.57828, 
    64.24458, 63.84927, 63.39538, 63.22643, 63.62318, 67.0251, 69.70273, 
    70.2049, 69.86025, 70.13414, 70.53278, 70.79231, 71.36761,
  91.99019, 92.29601, 92.64735, 93.07208, 93.47598, 93.75944, 94.08036, 
    94.35187, 92.82374, 92.98485, 93.15189, 93.83294, 93.88699, 93.75219, 
    94.38564, 94.23317, 93.54662, 93.70928, 94.16856, 94.05038,
  87.17807, 88.13142, 89.07693, 89.95754, 90.87383, 91.79653, 92.65139, 
    93.42416, 89.90855, 90.64588, 91.4202, 92.30596, 93.15186, 94.00761, 
    94.74245, 95.45621, 93.64816, 94.28283, 94.77159, 95.33623,
  85.98318, 87.58943, 89.21526, 90.60536, 91.84143, 93.05332, 94.14502, 
    95.07281, 90.72174, 91.58034, 92.57727, 93.43669, 94.46335, 95.25935, 
    95.93508, 96.69104, 95.19822, 95.96636, 96.59667, 97.01974,
  86.27484, 88.23713, 89.96051, 91.46679, 92.85941, 94.05687, 95.11847, 
    96.04095, 93.50178, 94.33504, 95.29518, 95.98656, 96.33752, 96.4943, 
    96.54282, 96.68465, 97.56662, 97.70418, 97.64644, 97.78993,
  84.76913, 87.29807, 89.51502, 91.14054, 92.5674, 93.68481, 94.33095, 
    94.8952, 94.01064, 94.24482, 94.66311, 95.02766, 95.36797, 95.57063, 
    95.89165, 95.48592, 97.79571, 97.19977, 96.49904, 95.97124,
  83.40446, 86.2171, 88.54231, 90.25722, 91.46258, 91.90891, 92.38571, 
    92.03294, 87.32184, 87.17188, 87.03313, 87.27244, 87.67892, 88.33023, 
    89.23311, 89.38163, 95.86903, 96.07491, 95.99859, 95.67516,
  88.73975, 87.60028, 87.66464, 88.93349, 89.56315, 89.47501, 88.89762, 
    88.81979, 80.98536, 79.7469, 76.43104, 76.72987, 77.56476, 81.31445, 
    82.82835, 82.1683, 89.16125, 91.48758, 93.44881, 94.06337,
  88.59106, 85.3774, 82.30107, 81.60769, 81.47722, 81.7335, 81.77341, 
    81.41296, 74.15842, 73.11501, 72.04942, 81.19814, 82.68713, 85.32762, 
    81.82372, 81.47345, 84.94654, 87.03708, 86.52367, 87.5546,
  81.48575, 80.28913, 78.38828, 76.62372, 75.64256, 75.48985, 75.38669, 
    75.02256, 72.86016, 73.68118, 74.48516, 75.47639, 77.76733, 80.44888, 
    82.00598, 82.48367, 81.67754, 81.75684, 87.41368, 91.02186,
  85.27977, 84.81836, 83.87429, 83.30049, 82.74548, 82.46806, 81.73237, 
    80.3901, 79.15118, 78.13171, 77.62334, 78.21085, 79.66831, 81.22745, 
    82.89187, 84.44139, 85.3705, 85.92397, 86.32735, 87.1496,
  88.64133, 88.61677, 88.10435, 87.60186, 87.9011, 88.53299, 88.78295, 
    88.30452, 86.95271, 84.76265, 82.37508, 81.55952, 81.96294, 83.07082, 
    84.14829, 84.58146, 84.42097, 84.13232, 84.02224, 84.81512,
  90.79475, 90.69728, 90.63476, 90.64536, 90.89552, 90.97123, 90.29098, 
    90.17594, 90.21941, 89.64416, 88.5708, 87.70496, 87.01369, 86.19238, 
    85.19343, 85.02781, 84.99041, 85.08275, 84.27575, 83.65764,
  92.73867, 92.4644, 91.92881, 91.58578, 90.7053, 88.67699, 85.5022, 83.7295, 
    83.73695, 84.6017, 84.79205, 85.27223, 86.34838, 87.16639, 87.43338, 
    87.02161, 87.59119, 88.01183, 87.11036, 85.60088,
  90.25692, 87.9325, 86.24883, 84.86899, 82.47671, 80.09042, 78.51436, 
    78.25417, 78.69518, 79.52922, 80.54766, 82.23596, 84.31653, 86.2239, 
    87.0758, 87.17768, 86.89486, 87.25323, 87.85658, 87.74698,
  88.03923, 83.48006, 79.07913, 77.03687, 75.91902, 75.81003, 76.54231, 
    77.39162, 78.22265, 79.38157, 81.27161, 83.12121, 84.76591, 85.25625, 
    84.52814, 84.25208, 84.4661, 85.13419, 86.44997, 87.83257,
  85.57114, 81.62355, 77.37597, 75.87283, 75.91644, 76.9922, 78.00246, 
    78.67866, 79.6945, 80.83163, 82.09543, 83.17196, 83.84315, 83.52836, 
    83.01657, 83.27694, 83.59528, 84.17583, 85.49647, 86.29888,
  81.90182, 79.94268, 78.98762, 79.36192, 79.44197, 79.40418, 78.99213, 
    78.62778, 78.54352, 79.06316, 79.62005, 80.52374, 81.2535, 81.94975, 
    81.99139, 82.06353, 81.36548, 80.97882, 81.28984, 81.41186,
  78.76537, 79.39391, 80.26613, 80.32736, 80.04203, 79.28844, 77.51565, 
    75.14468, 72.4982, 71.88822, 72.73312, 74.95419, 77.57262, 79.25433, 
    79.39274, 78.89417, 77.56009, 75.69604, 74.62907, 74.83327,
  76.06725, 76.28299, 75.37142, 75.3562, 76.31824, 76.1396, 72.65688, 
    66.7953, 63.30239, 61.70251, 61.48763, 63.67879, 68.22861, 71.73837, 
    72.27505, 71.72111, 70.25488, 68.54643, 67.82239, 67.84756,
  71.72768, 70.2263, 68.79956, 70.00876, 73.42229, 72.95086, 69.1363, 
    62.5623, 63.22075, 63.82442, 62.75166, 63.67667, 67.89378, 70.93182, 
    70.81177, 70.06979, 69.35578, 68.196, 67.06496, 66.68174,
  93.07325, 93.49728, 93.5911, 94.10221, 94.80148, 94.65248, 95.1761, 
    95.83871, 94.05556, 94.41294, 94.77554, 95.20275, 95.30827, 95.30733, 
    95.60662, 95.77581, 94.95175, 95.01777, 95.35828, 95.19642,
  85.55347, 86.76031, 88.06444, 89.27718, 90.58408, 91.78432, 92.95449, 
    94.01386, 90.60795, 91.40968, 92.08324, 92.74685, 93.62457, 94.58392, 
    95.35414, 96.31524, 94.88727, 95.5583, 96.07169, 96.68565,
  89.16733, 91.00497, 92.72155, 94.32832, 95.36557, 96.1729, 96.66209, 
    96.96385, 92.43015, 93.27235, 93.75489, 94.21878, 95.00962, 95.50878, 
    95.50539, 96.09323, 95.1252, 96.01401, 96.65579, 97.31917,
  88.10202, 90.30487, 92.26045, 93.71693, 94.82484, 95.62698, 96.40477, 
    97.06176, 95.41633, 96.30965, 96.52806, 97.19106, 96.96816, 96.78442, 
    97.13346, 98.29528, 99.13494, 99.05592, 98.95438, 98.70518,
  85.18156, 86.88393, 88.37735, 89.57432, 90.83894, 92.07703, 93.09739, 
    93.59739, 92.14561, 91.39977, 90.82958, 91.85632, 92.48899, 94.36236, 
    95.99239, 97.18658, 99.5212, 99.35587, 98.75349, 97.95295,
  82.52557, 84.40195, 86.09566, 87.8061, 88.92245, 89.67985, 89.88797, 
    89.88081, 85.36226, 85.41703, 86.05254, 86.86426, 87.83776, 89.01056, 
    89.7225, 90.75743, 96.69637, 97.01329, 96.99992, 96.28745,
  92.52042, 91.84008, 91.76089, 91.74084, 92.0473, 92.97919, 93.35713, 
    93.35458, 86.86846, 87.17076, 87.41853, 78.14487, 78.63598, 84.6556, 
    87.77859, 83.80342, 91.1165, 94.26971, 95.70324, 95.58753,
  88.04764, 85.22353, 83.19915, 83.37749, 83.65091, 86.27558, 88.88612, 
    89.15401, 83.51795, 83.44157, 83.25684, 81.31924, 82.44734, 89.5135, 
    90.55685, 91.77741, 92.1457, 92.06645, 87.49968, 87.96477,
  77.56745, 76.46099, 75.2754, 73.85542, 72.62728, 72.43127, 73.31264, 
    73.88206, 71.39237, 71.1645, 70.90585, 70.79633, 72.48635, 73.68194, 
    75.11298, 76.71381, 79.81185, 84.79149, 89.84075, 91.98466,
  82.25918, 82.3019, 82.22743, 82.13251, 81.87167, 81.42607, 80.49727, 
    79.47592, 78.70222, 78.05624, 77.46442, 76.60493, 75.84302, 74.66718, 
    72.53278, 70.59254, 69.52139, 69.87595, 71.11449, 72.41119,
  85.34775, 85.32586, 85.08144, 84.89854, 84.65031, 84.3327, 84.02703, 
    83.77882, 83.72484, 83.47941, 83.07838, 82.35089, 81.61643, 81.24581, 
    81.25786, 81.23319, 80.82311, 79.76589, 78.78503, 78.95351,
  86.6524, 86.81665, 87.36037, 88.23138, 88.58533, 88.39275, 87.50479, 
    87.54583, 88.07168, 87.78329, 87.00489, 86.423, 86.32674, 86.75478, 
    87.56242, 88.19028, 88.84011, 88.881, 87.08176, 85.42857,
  88.43851, 88.16961, 88.22265, 88.67272, 88.69275, 87.28993, 85.42874, 
    84.96664, 85.5114, 85.54277, 84.95732, 84.95036, 86.10343, 87.8328, 
    89.74329, 91.0747, 91.66318, 91.20206, 90.30211, 89.07913,
  86.92146, 84.9297, 83.63375, 83.47375, 82.81264, 81.34533, 80.73336, 
    81.22316, 82.40861, 83.25086, 83.87003, 85.00204, 86.93576, 89.24963, 
    91.62118, 92.87708, 92.48167, 92.00197, 92.15176, 92.11431,
  85.36416, 81.54705, 78.7467, 78.00748, 77.21777, 77.19073, 78.5243, 
    80.52879, 82.52884, 84.09219, 85.7934, 87.89032, 89.74417, 90.93546, 
    91.70303, 91.79339, 91.30603, 91.0872, 92.11804, 92.84982,
  83.0035, 79.60513, 76.12175, 75.9108, 76.57237, 77.94428, 80.42844, 
    82.28333, 83.43639, 84.80936, 86.2483, 87.30251, 87.75884, 87.86523, 
    87.35679, 86.86792, 86.46476, 86.7533, 88.12297, 88.53384,
  76.46925, 74.799, 74.44715, 76.24923, 78.01498, 79.64194, 80.56214, 
    80.79659, 80.96865, 81.36735, 82.17173, 82.7766, 82.89494, 83.27274, 
    82.83103, 81.72878, 80.26283, 79.60983, 79.8969, 80.46399,
  70.00018, 71.60336, 74.35414, 75.51313, 75.82394, 75.77158, 75.1762, 
    72.61008, 69.21627, 68.21412, 70.4205, 73.83517, 76.42325, 78.05372, 
    78.45387, 77.23768, 74.96582, 73.0297, 73.0284, 74.46644,
  67.5614, 69.07537, 69.36832, 68.95325, 69.20344, 68.61981, 65.69465, 
    61.36646, 59.10361, 58.07418, 58.54606, 59.86936, 62.00782, 64.63608, 
    67.13098, 68.25558, 68.96809, 69.95383, 71.67072, 73.26379,
  64.82347, 64.2474, 63.0896, 63.96076, 66.31025, 66.25845, 66.3396, 
    62.27503, 63.79876, 64.47713, 62.59331, 62.31839, 64.92087, 67.73288, 
    69.39334, 70.32552, 71.61484, 73.08654, 74.39008, 75.4177,
  92.93261, 93.28596, 93.35516, 93.81065, 94.4008, 94.2626, 95.00478, 
    95.33805, 93.75907, 94.01952, 94.36327, 94.54005, 94.62067, 95.06643, 
    95.15504, 95.3343, 94.40317, 95.00718, 94.85843, 95.46278,
  89.2488, 90.46349, 91.55478, 92.49122, 93.2949, 94.51505, 94.85549, 
    95.5313, 91.83494, 92.49745, 93.23412, 94.13586, 95.02124, 95.77672, 
    96.65413, 97.65862, 96.31862, 96.91248, 97.34779, 97.59739,
  88.84979, 90.39043, 91.61786, 92.34837, 93.091, 93.92904, 94.36205, 
    94.91117, 90.61463, 92.53421, 93.55143, 94.35366, 94.99853, 95.26904, 
    95.23031, 94.60111, 93.15002, 93.76711, 94.24011, 95.42512,
  88.00076, 89.81073, 91.43589, 92.40341, 93.12164, 94.54745, 95.95651, 
    97.07375, 95.5302, 96.94657, 97.55222, 97.74236, 98.30912, 98.8037, 
    99.23196, 99.43858, 99.14974, 98.4856, 97.92959, 97.06008,
  83.65375, 85.93964, 87.39673, 87.81788, 88.10492, 88.8746, 89.11161, 
    90.87273, 91.74634, 93.29364, 95.55354, 97.14935, 98.10722, 98.80382, 
    98.85238, 98.68919, 99.73923, 99.73515, 99.58132, 98.8223,
  83.88594, 85.94509, 87.54058, 87.7879, 86.61382, 85.75569, 85.07043, 
    84.46658, 80.43974, 81.42879, 82.93454, 84.88713, 87.06818, 89.01983, 
    90.42752, 91.7519, 97.49798, 97.60307, 97.43286, 96.69843,
  93.89215, 91.46745, 91.43824, 91.27988, 90.14403, 88.46506, 86.25547, 
    85.42378, 77.72659, 78.64615, 80.96256, 73.36821, 75.06286, 80.87564, 
    84.20646, 82.61795, 89.30502, 90.98363, 92.19983, 92.95459,
  92.85843, 92.02903, 90.42542, 88.70937, 87.62282, 87.77959, 88.6994, 
    89.92479, 85.03532, 85.93835, 89.86459, 84.70448, 85.58015, 90.13954, 
    93.68829, 89.39601, 93.48656, 90.56689, 90.10461, 90.41435,
  71.66845, 69.2281, 68.67253, 69.25183, 70.39448, 72.41589, 72.33153, 
    70.12503, 64.0294, 62.40294, 64.21779, 70.59789, 79.1424, 84.82327, 
    86.96243, 87.77832, 88.98431, 92.22002, 94.83298, 95.04214,
  75.87019, 74.48451, 73.25512, 71.869, 70.41154, 69.31786, 68.10583, 
    66.37885, 63.56535, 61.05518, 59.35479, 58.64373, 59.48762, 61.56434, 
    62.81791, 63.45252, 64.87772, 69.65203, 74.54262, 78.18998,
  80.84458, 80.2886, 79.36272, 77.88608, 77.17924, 76.78337, 76.4082, 
    76.08517, 75.45062, 73.7541, 71.44114, 69.32919, 67.72067, 66.83317, 
    67.05889, 67.13648, 66.69024, 66.17717, 66.2654, 67.27242,
  83.61317, 83.37717, 82.87971, 82.02672, 81.28289, 80.29768, 79.1301, 
    79.57936, 80.26623, 80.03362, 78.5396, 77.30704, 76.51955, 76.28717, 
    76.16076, 75.92508, 75.74409, 75.67424, 74.34867, 73.74129,
  84.28878, 84.2655, 84.23712, 84.36752, 83.73877, 81.52518, 78.74273, 
    77.30909, 77.07296, 76.72343, 76.09798, 76.40099, 77.90855, 80.28068, 
    81.97952, 82.94968, 82.84479, 81.75195, 80.55088, 79.98795,
  81.92359, 80.46687, 79.54182, 79.1226, 77.65541, 75.33714, 73.14993, 
    72.56432, 73.10941, 73.98235, 74.55755, 75.60131, 77.64203, 80.82716, 
    83.57835, 84.71386, 84.24144, 83.78573, 83.96893, 84.43049,
  81.71609, 78.00498, 73.94935, 71.65869, 69.87648, 68.29543, 67.47343, 
    68.49005, 70.63467, 72.86256, 74.79619, 77.19816, 79.90322, 82.27111, 
    83.73684, 84.35101, 84.19608, 83.83595, 84.31044, 85.50895,
  79.08899, 74.89923, 69.92703, 67.97023, 68.2564, 68.99601, 70.25818, 
    72.89051, 75.39928, 77.66824, 79.66955, 81.4472, 83.02357, 83.67107, 
    82.81256, 81.76521, 80.68292, 80.13757, 80.98457, 81.78413,
  75.06947, 72.29487, 71.19392, 72.46223, 73.98164, 75.59454, 76.85767, 
    78.11208, 78.74899, 79.36934, 79.85976, 80.16787, 80.6297, 80.75382, 
    79.75701, 78.33591, 76.34716, 74.78355, 74.10959, 73.46619,
  73.79073, 73.77792, 75.19384, 75.90292, 75.73274, 75.69099, 74.60593, 
    71.00009, 66.24703, 64.66167, 66.01723, 69.13483, 71.82573, 72.60545, 
    72.1272, 71.53222, 69.52093, 67.3181, 66.39082, 66.79581,
  72.1614, 72.62323, 71.60814, 69.65097, 69.27525, 68.68238, 65.89779, 
    61.80765, 59.66166, 58.06352, 57.18514, 57.14843, 58.06574, 59.12871, 
    60.26378, 61.70014, 63.32249, 65.08215, 66.4006, 68.04818,
  68.00304, 66.94242, 65.03395, 64.58286, 66.36487, 67.40664, 68.82734, 
    67.73259, 69.59308, 69.13939, 63.50457, 60.64816, 61.73365, 63.89784, 
    65.1422, 67.01325, 69.20506, 70.80837, 72.14099, 72.90908,
  92.94379, 93.19464, 93.59647, 93.84496, 94.34352, 94.68431, 94.97848, 
    95.25247, 94.08648, 94.39115, 94.70226, 94.85888, 95.16113, 95.47808, 
    95.62714, 95.73052, 94.95319, 94.96731, 95.28782, 95.58369,
  88.04927, 88.94574, 89.9554, 90.89842, 92.04098, 93.12331, 94.08083, 
    95.03392, 91.4965, 92.28862, 93.12339, 94.4173, 95.37405, 96.09498, 
    96.71964, 97.3345, 95.68687, 96.15768, 96.44368, 97.47002,
  86.06409, 87.4221, 88.825, 90.10931, 91.48856, 92.93662, 94.02368, 
    95.15239, 90.59263, 91.605, 92.72401, 93.5256, 94.46693, 95.62373, 
    96.57816, 97.42676, 96.94645, 98.00816, 98.97916, 99.48615,
  85.89458, 87.69509, 89.44688, 91.32862, 92.74494, 93.81109, 94.50379, 
    95.24732, 92.69022, 93.42876, 93.80505, 95.2047, 96.52749, 97.80505, 
    98.70736, 98.74198, 98.78911, 98.60011, 98.35406, 98.16121,
  83.83449, 85.68549, 87.0815, 87.85809, 88.66055, 90.01887, 90.15737, 
    91.09702, 90.63641, 91.15792, 91.80719, 92.06484, 92.69069, 93.93963, 
    95.05304, 95.93007, 98.84708, 99.0324, 98.86295, 97.72159,
  79.74782, 80.295, 81.24541, 82.21837, 83.37281, 84.94888, 86.21882, 
    86.9013, 82.76167, 82.94291, 83.73477, 84.72583, 85.77509, 87.13875, 
    88.86868, 90.6202, 97.1977, 98.21311, 98.35815, 97.47976,
  91.14445, 86.4252, 85.35013, 85.74377, 85.85769, 85.74764, 85.38925, 
    84.98888, 76.87714, 77.36929, 78.57041, 73.3685, 74.65974, 81.02254, 
    83.23959, 81.63152, 89.18919, 90.87275, 91.51616, 91.80245,
  94.76578, 94.00776, 94.22734, 94.26319, 94.3672, 94.34301, 94.8184, 
    95.53479, 90.81051, 92.13364, 93.93763, 90.70457, 91.42736, 94.84251, 
    95.13795, 88.1268, 94.11858, 95.64223, 89.63034, 90.43361,
  93.58887, 93.25885, 95.08118, 95.36527, 95.36735, 95.759, 96.21562, 
    96.33513, 94.6451, 95.14709, 96.15859, 96.6217, 96.47566, 96.37053, 
    95.98343, 95.39183, 96.44452, 97.46101, 97.54691, 96.77875,
  81.61471, 79.88601, 79.91869, 79.20672, 78.21996, 78.51543, 80.9189, 
    82.37521, 83.09317, 84.52047, 86.78239, 90.30573, 92.30305, 93.40726, 
    93.86562, 93.74401, 93.75922, 94.55804, 95.30284, 96.59673,
  73.47106, 72.93761, 72.08518, 70.08115, 67.60639, 66.40231, 66.12131, 
    66.36364, 67.05909, 67.32343, 67.57664, 67.95992, 69.06886, 69.82018, 
    69.58066, 69.45624, 69.67019, 69.18359, 67.51196, 68.67722,
  74.26826, 73.64842, 72.62998, 71.43037, 70.22768, 68.42289, 66.72757, 
    66.49924, 67.41609, 67.96642, 67.71156, 67.34223, 67.38374, 67.80056, 
    68.36843, 68.98007, 69.83394, 70.90362, 70.20972, 69.39864,
  76.41934, 76.6217, 76.28568, 75.69892, 74.37354, 71.94505, 69.55985, 
    68.6034, 69.02871, 69.40862, 69.19047, 69.26272, 70.11564, 72.1255, 
    75.06616, 77.49833, 78.91567, 79.18963, 77.83932, 75.70992,
  75.15558, 74.23958, 73.26668, 72.28411, 70.83237, 69.16295, 67.77824, 
    67.34296, 67.96751, 69.38661, 70.40996, 71.29166, 72.68134, 75.78059, 
    79.60584, 82.03364, 82.05332, 81.41279, 80.66559, 79.50532,
  73.3887, 70.67184, 67.84316, 66.75175, 66.07429, 65.65509, 65.54544, 
    65.90838, 67.83891, 70.59564, 73.19794, 75.2123, 76.80004, 79.24258, 
    81.37791, 82.05322, 81.15475, 80.13093, 80.20251, 80.93825,
  70.02901, 67.69292, 64.03734, 63.64212, 64.82023, 66.41711, 67.9389, 
    70.01379, 73.95454, 77.73234, 81.13875, 83.35262, 84.57528, 85.49307, 
    84.94127, 83.25422, 81.26731, 79.54998, 79.44937, 79.54614,
  64.93102, 63.83827, 64.61146, 68.51095, 71.55467, 73.60378, 75.5681, 
    77.57073, 79.86059, 82.04264, 84.09668, 85.53278, 86.18385, 86.49739, 
    85.29574, 83.43871, 80.5729, 77.87812, 76.13012, 74.51025,
  63.4729, 67.20568, 72.54038, 76.2365, 77.02151, 76.55251, 74.2457, 
    70.08839, 66.79724, 66.83519, 69.74707, 73.82656, 77.42665, 79.65483, 
    80.58582, 79.53799, 76.359, 71.94067, 68.88474, 67.98253,
  65.59491, 70.06881, 72.89611, 72.88049, 71.41888, 67.95296, 62.39409, 
    58.0667, 56.96686, 56.0612, 57.57288, 60.89142, 64.25356, 66.4799, 
    67.7486, 67.88627, 67.97484, 67.70634, 68.46278, 69.7133,
  63.73529, 65.25416, 65.93649, 66.41321, 65.46808, 63.71253, 63.43255, 
    63.86098, 65.41309, 65.2878, 61.07001, 61.94333, 65.64693, 67.32944, 
    67.28107, 68.97246, 72.1554, 74.44485, 75.33707, 75.00577,
  90.99626, 91.25625, 91.89591, 92.57214, 92.67012, 93.66508, 94.20377, 
    94.68235, 93.40678, 93.87612, 94.15051, 94.72164, 95.46111, 95.66187, 
    96.0202, 96.22688, 95.80862, 96.07925, 96.25059, 96.38721,
  85.27447, 86.65349, 88.18114, 89.55101, 90.93395, 92.23299, 93.22195, 
    94.39111, 91.17501, 92.08419, 92.90498, 93.89932, 94.86649, 95.82456, 
    96.62307, 97.22052, 95.74303, 96.80358, 97.36282, 97.9295,
  87.43353, 88.89176, 90.20712, 91.42925, 92.65008, 93.91302, 95.11971, 
    96.39597, 92.33887, 93.3653, 94.4939, 95.53975, 96.55833, 97.23904, 
    98.19843, 98.55145, 97.83423, 98.64576, 99.22348, 99.24442,
  88.87891, 90.94595, 92.74324, 94.29492, 95.18266, 95.61457, 96.30637, 
    96.62516, 94.25341, 94.9274, 95.75558, 96.87574, 97.6212, 98.25523, 
    98.8455, 99.24006, 99.53806, 99.51364, 99.29455, 98.64236,
  87.52349, 90.62015, 93.28596, 94.45826, 95.26169, 95.42973, 94.92532, 
    94.16565, 93.42338, 93.91051, 94.7049, 95.49426, 96.55215, 97.47273, 
    98.53236, 99.08961, 99.75945, 99.79984, 99.89714, 99.96413,
  83.01635, 84.30074, 85.23012, 85.86749, 86.59354, 87.74319, 88.60034, 
    88.86033, 84.04842, 83.77391, 84.46079, 85.64565, 87.33674, 89.14066, 
    90.71491, 92.15868, 98.11443, 98.45441, 98.26524, 97.56508,
  95.21119, 91.33134, 90.08892, 89.08617, 88.1017, 88.36624, 88.16536, 
    88.03094, 81.13039, 83.4175, 84.09683, 78.16368, 80.18185, 86.098, 
    88.1525, 84.1286, 89.34959, 90.75757, 91.80036, 92.31901,
  95.98233, 95.5732, 95.37262, 95.51505, 95.3912, 96.30369, 96.57922, 
    97.53994, 95.19373, 95.22156, 95.15201, 93.36585, 92.83157, 96.14072, 
    97.80115, 91.26502, 95.9001, 95.24105, 91.21841, 90.35344,
  99.53737, 99.37737, 99.07713, 98.96116, 98.59947, 97.95093, 96.86089, 
    96.63004, 94.3821, 94.9855, 96.0322, 96.90523, 97.61433, 97.20554, 
    97.39284, 98.42803, 98.9847, 99.1202, 98.58694, 97.34911,
  98.29868, 97.59079, 96.28345, 95.35509, 94.11423, 93.05286, 92.86745, 
    94.16303, 94.78882, 94.97315, 95.0816, 95.52547, 96.03916, 96.43701, 
    97.67091, 98.6911, 98.3847, 98.51966, 98.5044, 98.36401,
  92.45986, 93.66589, 93.75802, 94.69799, 94.83146, 93.12325, 90.70197, 
    90.97184, 91.99994, 92.49966, 92.19926, 92.06937, 92.41911, 92.76463, 
    93.68198, 93.94861, 93.90905, 93.84446, 91.64246, 88.29272,
  71.68362, 74.93998, 76.93916, 78.39185, 77.53773, 74.41798, 72.65017, 
    72.9995, 73.49395, 73.50494, 73.31072, 73.48769, 74.73997, 76.67753, 
    77.9475, 78.12567, 78.89252, 79.70976, 77.46385, 75.24524,
  74.38094, 76.05618, 77.38828, 78.93947, 79.45342, 78.35723, 76.55522, 
    75.69174, 75.81627, 76.04292, 76.25553, 76.696, 77.41821, 78.71535, 
    79.93114, 80.83792, 81.09782, 81.06504, 80.57716, 79.90873,
  74.95719, 74.49761, 74.41531, 75.10054, 75.26582, 74.6525, 74.2214, 
    74.91783, 76.63262, 78.19257, 79.29642, 80.38053, 81.6304, 83.05811, 
    84.94061, 86.70823, 86.40297, 85.61108, 85.29576, 85.33134,
  75.31238, 72.9622, 70.40456, 69.09753, 67.83889, 67.27892, 68.32871, 
    70.52743, 73.53821, 76.61526, 79.81371, 82.22334, 84.19176, 85.51209, 
    86.91376, 88.03082, 88.22648, 87.75847, 88.00953, 88.60606,
  75.0073, 71.60212, 66.29149, 62.97105, 62.18384, 64.02987, 67.40717, 
    70.53503, 74.8598, 79.28106, 82.85687, 85.26107, 86.86573, 88.31851, 
    88.76247, 88.37119, 87.7831, 87.4465, 87.89516, 87.91444,
  69.41142, 64.7308, 61.99051, 63.60659, 66.88065, 70.40561, 73.83842, 
    76.59113, 79.37697, 81.73637, 83.77877, 85.64483, 86.92168, 87.63211, 
    87.3689, 86.66803, 85.18652, 83.75054, 82.90009, 81.93539,
  66.62368, 67.67835, 70.9106, 74.07619, 75.49902, 75.9838, 74.59479, 
    70.56641, 67.32117, 66.26797, 68.0811, 72.30219, 77.13327, 79.18144, 
    80.25925, 79.95876, 76.98511, 72.45372, 69.3905, 68.31467,
  73.78598, 76.90626, 77.53636, 75.96872, 73.91189, 69.92731, 63.91581, 
    59.47733, 57.48041, 54.11458, 52.76872, 54.68633, 58.5851, 61.67231, 
    62.7364, 61.91265, 60.77544, 60.61396, 62.34473, 64.21873,
  74.83965, 75.02679, 72.79879, 70.60117, 68.49023, 66.29312, 65.0211, 
    66.45994, 66.37892, 63.37049, 57.1163, 56.72945, 60.70412, 63.65284, 
    62.87735, 61.38245, 62.53003, 64.85583, 68.46448, 70.6521,
  94.19295, 94.51764, 94.83413, 95.21857, 95.59444, 95.91167, 96.36088, 
    96.66115, 95.2778, 95.61436, 95.88277, 96.23495, 96.70492, 96.9987, 
    96.70753, 97.18075, 96.62346, 97.06754, 97.07039, 96.84184,
  89.30978, 90.28778, 91.21302, 92.08656, 93.0288, 93.97791, 94.84388, 
    95.53498, 91.72358, 92.37656, 93.18641, 93.56998, 94.46183, 95.47736, 
    96.76683, 97.48086, 96.18582, 96.86652, 97.53548, 97.46899,
  87.37196, 88.92744, 90.42233, 91.6684, 92.73918, 93.38722, 94.46523, 
    95.30933, 90.80748, 92.15386, 93.3385, 94.72986, 95.78529, 96.05679, 
    96.74356, 97.43968, 97.2037, 97.652, 98.12968, 98.73502,
  87.6966, 89.62521, 91.50441, 92.91175, 93.96711, 95.26143, 96.40824, 
    97.10127, 95.01966, 95.24596, 95.63797, 96.42078, 97.08805, 98.07513, 
    99.01602, 99.56732, 99.71205, 99.49722, 99.02661, 98.24929,
  86.8343, 88.76755, 89.46332, 90.54125, 91.52932, 92.16376, 92.0174, 
    93.15366, 93.85455, 94.58593, 94.65598, 95.17631, 96.02085, 97.03032, 
    97.66964, 98.1329, 99.49753, 99.80218, 99.85336, 99.80305,
  80.98493, 81.18821, 82.74544, 83.95581, 84.68581, 85.36117, 85.79142, 
    86.59299, 83.16241, 84.04737, 85.14357, 86.30415, 87.50468, 89.16687, 
    90.8682, 92.27048, 97.42408, 98.09206, 98.42406, 98.0501,
  91.66521, 87.61363, 86.17207, 86.33651, 86.31835, 85.99666, 86.14391, 
    85.84721, 78.35093, 78.49154, 79.88809, 75.47124, 78.33195, 86.6847, 
    87.93015, 86.79314, 92.75163, 93.81, 94.4985, 94.38663,
  96.93368, 96.30988, 96.22165, 96.84893, 97.57732, 97.15742, 97.18052, 
    96.49612, 94.38546, 94.72186, 96.27824, 95.53788, 95.47644, 97.16564, 
    98.06435, 89.56399, 95.49038, 94.83575, 91.71381, 92.08071,
  97.0528, 97.30752, 96.97052, 96.19128, 97.10697, 97.82839, 97.87937, 
    97.14817, 95.3354, 96.7373, 97.37254, 98.16196, 98.59366, 99.06174, 
    99.13651, 99.40726, 99.55504, 99.77026, 99.40911, 98.89939,
  94.97549, 96.77702, 97.41358, 97.41988, 97.23911, 97.04185, 96.92985, 
    95.49656, 93.25801, 93.00709, 93.76648, 94.2645, 95.68218, 96.21618, 
    96.50294, 97.09788, 97.3086, 98.33789, 98.85184, 98.88365,
  94.27692, 95.35107, 97.2251, 97.86195, 97.77716, 97.73415, 97.40862, 
    96.48288, 95.2018, 96.66145, 97.33264, 97.21115, 97.10863, 97.34924, 
    97.3121, 96.66038, 95.60918, 95.33842, 94.24186, 92.50967,
  91.47499, 92.33476, 93.00029, 94.17915, 93.85282, 85.12591, 72.89086, 
    71.02183, 74.01675, 76.01976, 76.07388, 75.75114, 76.40945, 80.54135, 
    87.79263, 90.74916, 92.47885, 93.89842, 89.32902, 81.7963,
  71.38752, 72.24569, 72.69078, 73.22079, 72.78973, 70.34103, 67.9206, 
    67.07028, 67.18874, 67.80492, 68.15817, 68.14363, 68.7894, 70.19366, 
    72.12502, 73.64125, 74.11829, 74.61341, 73.10235, 69.74648,
  70.54379, 70.09124, 70.22389, 71.91786, 72.90658, 73.09746, 72.77913, 
    72.80836, 73.9738, 75.53783, 76.20168, 76.72182, 77.4728, 78.03043, 
    78.77598, 79.71165, 79.1304, 78.47903, 77.79527, 76.26522,
  72.54208, 71.82574, 71.03272, 71.15619, 70.11339, 69.45035, 69.3802, 
    70.54711, 73.1226, 75.49863, 77.49395, 79.46597, 80.80301, 81.27815, 
    81.46027, 81.9041, 81.32973, 80.07281, 79.07342, 78.62608,
  71.4409, 70.53636, 67.30802, 65.39652, 64.84406, 65.70407, 68.063, 
    71.33327, 76.08868, 80.585, 84.03281, 85.94774, 86.58956, 86.63538, 
    85.97544, 84.45186, 81.54161, 78.50562, 77.39528, 76.97617,
  66.42821, 63.1954, 61.25183, 63.47744, 66.69307, 70.7377, 75.00713, 
    79.10089, 83.27927, 85.99637, 87.88502, 89.03252, 89.52077, 88.86276, 
    86.90957, 83.91634, 79.01649, 74.59162, 71.52484, 69.7934,
  60.13446, 62.85339, 67.75481, 72.25069, 75.71808, 78.21542, 78.47874, 
    76.26804, 73.4269, 71.96439, 73.25713, 76.66979, 80.07168, 81.30844, 
    80.63612, 77.9703, 72.06354, 65.94221, 62.62874, 61.25689,
  66.21132, 70.73206, 73.82254, 75.29621, 74.55597, 71.12618, 65.87658, 
    62.08369, 60.66447, 58.24749, 57.32602, 58.96198, 62.58973, 65.00629, 
    65.35915, 64.06774, 61.24484, 59.27686, 59.26825, 60.20398,
  68.73228, 70.32368, 70.90421, 70.77377, 68.29355, 64.97314, 63.21965, 
    63.76423, 66.17312, 64.82809, 59.11375, 59.34901, 64.39133, 67.8831, 
    66.94431, 65.66779, 64.84155, 64.37527, 64.77981, 65.15578,
  93.51248, 93.77986, 94.2194, 94.44169, 94.60114, 94.94878, 95.26913, 
    95.51363, 93.96811, 94.47356, 94.4088, 94.82061, 95.21985, 95.09193, 
    95.46581, 95.79934, 94.58129, 94.6806, 95.64635, 95.46514,
  85.53738, 87.03603, 88.59386, 90.07538, 91.45131, 92.67375, 93.78709, 
    94.71454, 91.6599, 92.54829, 93.50476, 94.34512, 95.2797, 95.91132, 
    96.59088, 97.39109, 96.63418, 96.96376, 96.98259, 97.16312,
  85.23771, 87.6843, 89.96255, 91.80358, 93.14434, 93.92175, 94.9016, 
    95.69683, 91.17004, 91.12202, 91.34238, 92.72179, 93.87966, 94.56243, 
    94.99118, 95.66899, 95.20592, 95.97505, 97.16917, 98.33385,
  87.79712, 89.98769, 91.97586, 93.24567, 94.22997, 95.48856, 96.45098, 
    96.99919, 95.24645, 95.97117, 96.86954, 97.77989, 98.44939, 98.74747, 
    99.09893, 99.44555, 99.55146, 99.4364, 99.12006, 98.61757,
  80.99118, 83.4847, 85.91704, 87.81411, 89.56752, 91.4834, 92.99966, 
    94.31182, 94.49595, 94.85894, 95.22187, 95.59814, 95.92651, 95.83332, 
    95.29397, 96.10369, 98.29241, 98.07743, 98.52029, 99.28881,
  80.04578, 82.61535, 84.76769, 86.25637, 87.45481, 88.42133, 88.91893, 
    88.81651, 84.18646, 84.1218, 84.9787, 86.03481, 87.12576, 88.12206, 
    89.10474, 89.97378, 95.69219, 96.80936, 97.84075, 97.47741,
  92.55618, 90.2897, 89.98019, 90.53651, 90.85149, 90.6901, 90.1814, 
    89.48147, 81.61734, 81.71169, 82.05006, 76.23808, 77.55069, 84.22401, 
    84.77674, 80.58569, 86.95667, 88.98992, 90.29689, 90.59538,
  97.98399, 98.03358, 98.1911, 98.51582, 99.17842, 99.31967, 98.98422, 
    98.79011, 94.85764, 95.63545, 94.12568, 94.51499, 94.6152, 97.50035, 
    97.65218, 89.71871, 94.38531, 92.25273, 85.66553, 86.21886,
  98.51627, 99.18169, 99.3055, 99.09796, 98.98017, 98.71434, 98.35857, 
    98.24113, 97.30846, 97.62593, 97.91573, 98.17841, 98.42879, 98.47256, 
    98.75642, 99.04606, 98.74485, 99.00974, 98.91488, 98.4099,
  97.37083, 97.22188, 97.06409, 97.12318, 97.03062, 96.69138, 96.39138, 
    96.07223, 96.31979, 97.44938, 98.3774, 98.46991, 98.21931, 98.00174, 
    98.17706, 98.46072, 98.31724, 98.82293, 99.10559, 99.3125,
  96.13039, 96.10419, 95.88728, 95.99425, 95.81258, 95.3777, 94.96558, 
    94.95728, 95.5175, 96.13953, 96.59737, 96.79588, 96.85063, 96.7679, 
    96.69569, 96.61954, 95.72032, 96.05701, 96.3499, 96.58568,
  92.37275, 92.0697, 91.19598, 91.24213, 92.65855, 92.00672, 86.31123, 
    83.2442, 82.56106, 82.78432, 83.47523, 84.18024, 87.02102, 90.9268, 
    92.69891, 93.31573, 92.80495, 93.54334, 94.04441, 90.75733,
  78.06488, 79.15591, 79.62674, 79.54352, 78.56039, 75.10004, 70.67941, 
    68.62946, 68.30299, 68.06812, 67.51235, 67.29737, 68.41395, 70.62189, 
    72.81313, 74.26956, 74.89629, 76.72488, 77.01946, 74.42144,
  77.73622, 76.95366, 76.21229, 75.8689, 74.95994, 73.47634, 71.6442, 
    70.10614, 69.49809, 69.94774, 70.77177, 72.36104, 74.88303, 77.35417, 
    78.69822, 79.00974, 77.97067, 77.49902, 77.6906, 77.42421,
  81.04718, 79.38941, 77.43924, 76.16879, 74.29528, 72.15816, 70.58189, 
    69.76585, 70.41129, 72.47678, 75.36807, 78.48029, 81.19725, 82.61316, 
    82.82358, 82.99673, 82.93633, 82.98636, 83.24992, 84.21691,
  81.21257, 79.08103, 74.41717, 69.6515, 66.76323, 65.78361, 65.79103, 
    67.16759, 70.85918, 75.40105, 79.51749, 82.49249, 84.2086, 85.17521, 
    85.52007, 85.48971, 84.13799, 82.3965, 82.18932, 82.72845,
  75.58995, 70.05966, 63.76106, 61.51537, 62.23551, 63.76125, 65.9638, 
    69.13084, 72.53968, 76.13222, 79.74849, 82.73069, 84.60073, 85.36042, 
    84.96481, 83.55095, 80.40121, 77.42368, 75.46912, 73.75533,
  64.26098, 63.85443, 65.89986, 66.74401, 69.31903, 71.32278, 71.76369, 
    69.42471, 66.94117, 66.36002, 67.94485, 70.98315, 74.31165, 75.76672, 
    75.97987, 75.3274, 71.8425, 67.35387, 64.4713, 62.91702,
  68.83983, 70.90859, 71.36927, 71.55132, 71.21906, 68.89108, 65.58945, 
    63.10664, 61.38224, 58.71861, 57.38202, 58.77856, 61.49718, 63.77268, 
    65.59793, 66.10002, 65.10695, 63.78395, 62.94027, 63.05755,
  70.32998, 69.08137, 68.34586, 68.5285, 67.32476, 65.13901, 65.29192, 
    68.19952, 69.3458, 67.10061, 61.71188, 61.19221, 66.91853, 70.15424, 
    69.9238, 69.85007, 70.6242, 71.39331, 72.15957, 72.92717,
  90.41528, 90.90757, 91.2857, 91.78419, 92.13621, 92.52325, 92.86205, 
    93.12434, 91.66921, 92.18816, 92.52222, 92.79023, 93.17219, 93.42892, 
    93.89518, 94.23495, 93.4203, 93.52059, 93.70576, 94.05851,
  83.60858, 85.06452, 86.78461, 88.49007, 90.23019, 91.74763, 92.89125, 
    93.50168, 89.54099, 90.36035, 91.22127, 92.23608, 93.61193, 94.7267, 
    96.0038, 97.30542, 96.4469, 97.16927, 97.80681, 98.41525,
  83.11462, 85.37621, 87.50964, 89.64908, 91.25517, 92.07388, 92.94077, 
    93.66452, 89.21827, 89.45448, 90.17455, 92.08837, 93.19067, 94.62781, 
    95.76443, 96.51012, 96.05116, 96.68564, 97.50332, 98.30514,
  83.12463, 85.43916, 87.63168, 89.78548, 91.52615, 93.0627, 93.43797, 
    93.71944, 91.65083, 92.24783, 92.98074, 93.94497, 95.31674, 97.18475, 
    98.49461, 99.07525, 99.40901, 99.26551, 98.84558, 98.5359,
  80.2645, 81.91017, 83.37834, 84.73576, 85.01307, 85.21658, 85.53509, 
    86.33228, 86.37237, 87.95909, 89.92072, 91.8527, 93.64651, 95.0559, 
    96.4692, 97.33475, 99.12011, 99.41328, 99.60923, 99.35943,
  78.34957, 80.17643, 81.44513, 82.38741, 82.87919, 83.87804, 84.84511, 
    85.885, 82.40596, 82.83447, 83.44231, 84.62518, 85.566, 86.74519, 
    87.6605, 88.65749, 95.63538, 96.88885, 97.6991, 97.64062,
  91.8741, 89.66988, 89.32726, 89.25298, 89.12035, 89.39587, 89.23623, 
    89.95338, 82.81219, 83.46056, 85.60861, 76.79867, 78.55482, 86.48648, 
    88.5061, 85.38651, 91.81134, 93.11494, 94.1008, 94.31271,
  98.04394, 97.74216, 97.52959, 97.09235, 97.63771, 98.11301, 98.15636, 
    98.4482, 92.79355, 92.26116, 92.68295, 90.21172, 91.60065, 95.76173, 
    98.11726, 89.72677, 95.75099, 94.60648, 90.98551, 90.27503,
  97.70024, 97.72186, 97.43939, 97.39436, 96.85804, 96.59498, 96.04434, 
    94.16602, 90.44881, 90.88785, 92.8157, 94.42545, 95.42844, 95.88759, 
    95.79005, 96.42085, 97.16113, 98.58304, 98.33988, 98.19882,
  97.37814, 97.07377, 96.36613, 95.59668, 94.64588, 94.03108, 93.75379, 
    93.45353, 93.40286, 93.15197, 92.77137, 93.72333, 95.38643, 96.28882, 
    96.44494, 96.53462, 96.84122, 97.15372, 97.45715, 97.75092,
  96.7508, 96.69188, 96.39793, 96.37955, 96.59979, 96.63687, 95.69971, 
    95.06281, 94.87547, 94.70735, 94.37086, 93.99979, 93.89398, 94.07125, 
    94.34059, 94.58717, 95.25436, 95.2407, 95.55763, 95.71384,
  93.69402, 93.74519, 94.3308, 94.77013, 94.34531, 93.74538, 91.77161, 
    88.63348, 87.50249, 86.10595, 84.11406, 83.15276, 82.67438, 85.55404, 
    88.05633, 90.09569, 91.16019, 91.27743, 91.4013, 91.43288,
  82.10684, 82.23656, 81.64877, 81.06386, 80.07531, 77.19688, 71.52119, 
    67.48171, 67.08885, 67.72493, 68.02104, 68.74521, 70.21001, 72.76281, 
    75.46922, 77.38937, 78.76537, 79.89774, 81.55592, 80.89756,
  71.43602, 69.91088, 68.59511, 67.80733, 66.56128, 65.13577, 64.22041, 
    63.91716, 64.72094, 66.16068, 67.59854, 69.81393, 73.02245, 76.71758, 
    79.89941, 81.22356, 80.64238, 79.97198, 80.11705, 80.19773,
  73.55518, 70.82188, 68.10629, 66.43543, 64.44555, 63.11603, 63.17065, 
    64.1178, 66.30262, 69.24272, 72.64149, 76.40441, 79.72997, 82.15014, 
    83.19288, 83.47129, 83.43078, 83.88261, 84.5869, 85.39837,
  75.80796, 73.52658, 68.39201, 64.43924, 62.52713, 62.50118, 63.61297, 
    65.2522, 68.78353, 73.56409, 78.13705, 81.51473, 83.66412, 85.00379, 
    85.5891, 86.44411, 86.55976, 85.61225, 84.8504, 84.69051,
  71.30258, 66.69501, 62.08947, 61.57819, 62.84948, 64.59985, 66.54852, 
    68.887, 72.21695, 75.72128, 79.51714, 82.57623, 84.26987, 85.15051, 
    85.6331, 85.97474, 84.25445, 81.56079, 79.14803, 77.35355,
  62.97787, 63.61786, 67.24549, 69.73798, 71.23629, 72.46666, 72.99273, 
    70.84603, 68.28699, 67.86405, 70.26612, 73.54825, 76.36868, 78.13901, 
    79.00428, 78.72938, 75.11478, 70.08523, 66.95837, 65.85214,
  69.83939, 73.27724, 75.57932, 75.89419, 74.26587, 71.04425, 65.81826, 
    61.37852, 59.3793, 57.52807, 57.31192, 58.97566, 60.77186, 61.26305, 
    61.43164, 61.04893, 59.81348, 59.2662, 60.26337, 62.04465,
  72.89191, 72.77204, 72.19234, 70.51865, 67.49791, 65.5778, 64.77446, 
    63.62363, 64.87605, 63.39087, 59.4991, 58.32731, 61.18675, 62.15475, 
    61.50454, 61.41556, 62.22366, 64.04356, 66.53925, 68.97784,
  88.73393, 89.09306, 89.40646, 89.74352, 90.10521, 90.4968, 90.85628, 
    91.21909, 89.79095, 90.05299, 90.33064, 90.55548, 90.82059, 91.18579, 
    91.48916, 91.77986, 91.1551, 91.59414, 91.82942, 92.09741,
  81.30318, 82.36691, 83.5713, 84.92404, 86.32867, 87.7026, 89.1825, 90.5865, 
    87.59962, 88.7904, 89.65603, 90.37893, 91.16689, 92.05873, 93.0955, 
    94.15909, 92.66403, 93.78323, 94.75829, 95.62593,
  79.99127, 81.87746, 83.82252, 85.79079, 87.6862, 89.26919, 90.58695, 
    91.72974, 87.53243, 88.59083, 89.64082, 91.30486, 92.45798, 93.92944, 
    95.22604, 96.35035, 95.17547, 96.02132, 96.61123, 97.14442,
  80.7509, 83.46567, 86.17308, 88.56691, 90.70527, 92.5304, 93.59359, 
    94.22161, 91.98536, 92.99194, 94.20657, 95.53143, 96.72235, 97.48035, 
    97.83039, 98.01574, 98.62408, 98.59712, 98.20957, 98.0063,
  79.87002, 82.98624, 86.32561, 88.96359, 91.09431, 92.76335, 94.10354, 
    95.02315, 94.11189, 94.57732, 95.10331, 95.73466, 96.17744, 96.63283, 
    96.98975, 97.00783, 99.50397, 99.42043, 98.9466, 98.44539,
  80.76653, 83.46317, 85.6234, 87.95914, 89.8281, 91.05721, 91.61433, 
    91.82983, 87.54727, 87.58215, 87.9446, 88.55104, 89.40746, 90.48811, 
    91.61696, 92.57008, 97.87291, 98.07755, 97.98794, 97.40128,
  92.12874, 90.73962, 89.96543, 90.07652, 90.81475, 91.7746, 91.3423, 
    90.58308, 82.67265, 82.64446, 83.14261, 80.46693, 82.15479, 87.15137, 
    88.2571, 88.41931, 93.80453, 94.1982, 94.67073, 94.84233,
  95.60722, 94.99995, 94.17903, 93.751, 94.53782, 95.31149, 94.45164, 
    93.4188, 89.49586, 90.96862, 90.48697, 89.41054, 90.21236, 93.11912, 
    94.32756, 85.17836, 92.94205, 94.14449, 93.66626, 94.62081,
  95.55025, 95.5012, 95.12073, 94.37926, 94.15147, 93.43069, 92.50136, 
    92.74953, 91.78094, 93.2272, 93.135, 93.08343, 93.19742, 93.49413, 
    93.69791, 94.52171, 95.17285, 96.70741, 96.20411, 95.4704,
  94.656, 94.91176, 94.57431, 94.28602, 94.32684, 93.91409, 93.35975, 
    93.64709, 94.96495, 95.53642, 95.67834, 94.9754, 94.55679, 94.51383, 
    94.64596, 95.15974, 95.80762, 96.42763, 97.06981, 97.13276,
  94.97238, 94.80089, 94.47847, 94.47744, 94.44065, 94.13998, 93.61167, 
    92.93638, 93.15556, 93.89497, 94.71803, 94.39438, 93.83284, 93.89143, 
    93.74859, 94.02999, 94.48288, 94.21182, 94.31651, 94.17271,
  95.01912, 94.37193, 93.39437, 92.51048, 91.6839, 91.31615, 90.41712, 
    88.52367, 87.0819, 86.7802, 85.22184, 84.53474, 83.8605, 85.32542, 
    88.43973, 90.10593, 91.03016, 91.36336, 90.9447, 88.88686,
  88.83278, 86.61138, 85.06744, 83.56402, 81.25322, 77.45995, 71.46197, 
    66.5329, 64.83114, 64.50209, 64.1516, 64.76105, 66.90791, 70.81298, 
    75.2915, 77.89698, 79.15145, 79.62096, 79.87476, 79.49873,
  75.82814, 73.42361, 70.45572, 67.50496, 65.00971, 62.69215, 61.02328, 
    60.19524, 60.30513, 61.33287, 62.28439, 64.29026, 67.85814, 72.18125, 
    75.72052, 77.40501, 77.07944, 76.7822, 77.94156, 79.1611,
  76.32951, 73.50486, 69.6469, 66.0994, 62.45071, 59.59464, 58.27341, 
    58.42602, 59.44012, 61.87917, 64.78407, 68.48234, 72.41747, 75.50575, 
    77.24635, 77.49911, 77.16858, 77.20598, 78.36996, 80.1302,
  75.25082, 72.26967, 66.60489, 61.5107, 59.03014, 58.21657, 58.53315, 
    59.68136, 61.81092, 65.70576, 70.29401, 74.11465, 77.24475, 79.78107, 
    80.87707, 81.42825, 81.46172, 79.82925, 78.57266, 78.46312,
  71.47084, 66.25894, 61.0493, 59.98388, 60.7786, 62.13651, 63.57935, 
    65.18848, 67.10448, 69.95617, 73.33553, 76.27291, 78.66802, 80.70388, 
    82.30074, 83.60021, 82.20904, 77.77615, 73.84319, 71.76165,
  65.513, 64.47814, 67.05786, 68.50641, 70.1423, 71.89009, 72.61584, 
    69.43517, 65.12684, 64.39009, 66.54393, 69.84029, 74.01795, 77.27647, 
    79.51016, 79.54911, 75.77275, 69.30941, 64.84113, 63.24535,
  69.29553, 72.04801, 73.14484, 74.103, 73.72565, 71.20961, 65.54259, 
    60.00912, 55.53934, 53.28321, 53.3075, 55.69744, 59.52451, 63.17377, 
    66.23524, 67.1547, 65.95627, 64.36916, 63.92494, 64.55632,
  69.78914, 70.25249, 69.83482, 68.99891, 67.24076, 64.89074, 62.21782, 
    59.61015, 57.71795, 58.74483, 57.66247, 58.20327, 63.76088, 68.42136, 
    69.93115, 70.18614, 70.66887, 71.25742, 72.65355, 73.80934,
  88.38089, 88.73958, 89.11292, 89.43459, 89.78239, 90.15271, 90.50674, 
    90.88435, 89.27608, 89.54887, 89.8127, 90.11781, 90.31442, 90.62109, 
    90.81635, 91.1181, 90.37646, 90.4733, 90.71027, 90.74872,
  83.81244, 84.60059, 85.42902, 86.29432, 87.22014, 88.10642, 89.00329, 
    89.92122, 86.422, 87.27882, 88.1835, 88.96567, 89.78199, 90.63076, 
    91.57196, 92.44102, 90.68935, 91.3783, 92.04385, 92.73872,
  84.59193, 85.91069, 87.25675, 88.56311, 89.84476, 91.16595, 92.22168, 
    93.11965, 88.55827, 89.32095, 89.95499, 91.01475, 91.80087, 93.17109, 
    94.19267, 95.23058, 93.77059, 94.78114, 95.50777, 96.10487,
  85.56222, 87.49435, 89.28156, 90.83591, 92.3578, 93.65998, 94.57954, 
    95.45421, 92.81277, 93.38946, 93.82822, 94.26481, 94.72793, 95.33896, 
    95.81667, 96.30344, 97.29507, 97.30553, 97.19147, 97.12607,
  83.93439, 86.30239, 88.67644, 90.03889, 91.46249, 92.69587, 93.89952, 
    94.76527, 93.31333, 93.65929, 94.11357, 94.57063, 94.97847, 95.35831, 
    95.62093, 95.62465, 98.88004, 98.32402, 97.65939, 97.1028,
  82.54654, 85.26759, 87.32928, 88.87653, 90.08569, 90.63774, 91.23608, 
    91.66594, 87.41085, 87.83167, 88.7002, 89.75012, 90.73042, 91.64233, 
    92.40926, 93.37399, 98.65119, 98.5732, 98.18204, 97.52835,
  89.05071, 87.5925, 87.22859, 87.76056, 87.94604, 87.98019, 87.84013, 
    87.86852, 80.68434, 81.41273, 80.04623, 78.77972, 80.20045, 85.21616, 
    87.2953, 86.99444, 93.81437, 95.66595, 96.60863, 96.61929,
  90.37669, 91.02873, 91.27276, 91.56992, 91.56002, 91.18902, 90.9306, 
    90.69083, 86.26799, 86.01791, 82.16679, 83.24733, 84.23017, 88.93907, 
    92.20876, 83.51116, 89.16639, 92.30609, 91.9535, 94.19427,
  94.34652, 93.84478, 93.45161, 92.78756, 92.18559, 92.22164, 92.07063, 
    91.80862, 90.26094, 90.30153, 90.15939, 90.13844, 90.15646, 90.17203, 
    90.58335, 91.36133, 91.61637, 92.30571, 89.73852, 91.28978,
  96.73876, 96.38221, 95.9465, 94.85227, 93.909, 94.15883, 94.24763, 94.1897, 
    94.36102, 94.36282, 94.72205, 95.19411, 95.56963, 95.83561, 95.54597, 
    95.18438, 94.79053, 94.77996, 94.89502, 94.67316,
  95.44107, 95.63583, 95.66611, 95.1993, 94.22476, 94.40013, 94.79672, 
    95.36417, 96.08137, 96.41478, 96.48111, 96.12822, 95.99815, 96.48031, 
    96.23035, 96.10214, 95.57073, 95.44093, 94.98611, 94.75494,
  94.58598, 94.22112, 94.01154, 93.5696, 93.2723, 93.19897, 93.06255, 
    93.30874, 93.56513, 94.09024, 93.98666, 93.11509, 92.79926, 93.2181, 
    92.91521, 91.2878, 89.1066, 88.42892, 88.9345, 89.44263,
  92.75383, 91.98829, 90.58488, 89.62826, 88.47351, 85.89405, 82.47783, 
    80.49537, 79.39468, 77.99252, 76.50561, 76.45111, 78.28342, 81.02877, 
    83.55005, 84.48124, 84.59111, 85.1638, 86.18997, 86.80143,
  87.18379, 85.11624, 83.00953, 81.01562, 78.51731, 75.96429, 73.94781, 
    73.02708, 72.57465, 72.70415, 72.54212, 73.56361, 76.23782, 79.8047, 
    83.45802, 85.66119, 84.95119, 84.11485, 84.48538, 85.48387,
  87.1711, 84.16714, 80.01141, 76.32097, 72.65127, 69.75251, 68.56142, 
    68.23073, 68.26509, 69.10501, 70.90445, 73.44359, 76.66566, 79.74068, 
    82.32116, 83.86383, 83.32977, 82.38044, 83.09478, 85.09015,
  84.61023, 81.65151, 75.42706, 69.82507, 66.77296, 65.87753, 66.28108, 
    66.76443, 67.68835, 70.01642, 73.58195, 76.80556, 79.72779, 82.4463, 
    83.8488, 84.58154, 84.59566, 84.18756, 84.39393, 85.03338,
  79.68078, 75.17267, 69.04591, 67.55859, 68.13799, 68.79106, 69.07079, 
    69.39734, 70.31207, 72.27117, 74.7827, 77.3352, 79.70182, 81.80283, 
    82.95721, 83.60415, 83.1889, 81.96506, 80.19306, 78.10758,
  74.67362, 73.13733, 75.00191, 76.24243, 76.61693, 76.95782, 76.16199, 
    71.98969, 66.73979, 64.95311, 65.60272, 68.00574, 71.467, 74.36266, 
    76.25246, 76.75824, 73.96067, 69.75085, 66.79626, 65.43329,
  76.24976, 79.17164, 80.34796, 79.72572, 78.23902, 75.43619, 69.32655, 
    63.22482, 58.38475, 55.09309, 53.2612, 53.39599, 56.02224, 60.02954, 
    63.22612, 63.61857, 62.03452, 61.08965, 61.65327, 63.27081,
  75.27863, 75.36452, 74.26022, 73.04491, 71.26729, 68.45264, 65.17984, 
    62.36742, 62.71459, 60.83821, 56.34679, 54.55258, 58.32462, 62.31729, 
    64.06691, 63.74149, 63.79243, 64.9463, 67.36145, 70.35558,
  93.80733, 94.14867, 94.19357, 94.42138, 94.76548, 95.01586, 95.27175, 
    95.59641, 94.03018, 94.27721, 94.52475, 94.7265, 94.96246, 95.25582, 
    95.38172, 95.68968, 94.9475, 95.17612, 95.50465, 95.62811,
  84.60175, 85.52145, 86.67049, 87.7821, 88.68864, 89.88702, 90.79393, 
    91.74097, 88.32588, 89.16046, 89.88966, 90.74709, 91.47072, 92.19707, 
    92.87318, 93.55532, 91.63522, 92.18565, 92.47121, 92.98089,
  80.72478, 82.27682, 83.78984, 85.331, 86.96612, 88.4213, 89.80935, 
    90.81035, 86.60482, 87.64497, 88.51456, 89.2051, 90.10258, 90.82879, 
    91.44873, 92.2084, 90.16816, 90.85198, 91.26053, 91.73514,
  81.79185, 84.00179, 86.02912, 88.16181, 89.61056, 91.23441, 92.25012, 
    93.2299, 90.0988, 90.56508, 90.73689, 91.19297, 91.64268, 91.83379, 
    92.19187, 92.55071, 93.29836, 93.30566, 93.24217, 92.72644,
  81.58612, 84.54649, 87.05977, 89.39727, 90.78487, 91.90458, 92.62467, 
    92.80562, 91.029, 90.96974, 90.97515, 91.45186, 91.59333, 92.34634, 
    92.78953, 92.6869, 97.08359, 96.80997, 95.95485, 95.0303,
  82.27006, 85.27258, 87.88934, 89.74826, 90.88569, 91.37885, 91.56381, 
    91.60824, 87.02969, 87.10664, 87.26767, 88.03686, 89.23933, 90.11772, 
    91.81406, 92.90449, 98.52608, 98.36727, 97.89836, 97.13451,
  88.1868, 85.896, 85.76717, 86.52961, 86.75871, 86.61211, 86.06303, 
    85.63349, 77.71236, 77.01421, 75.14199, 76.18558, 77.37888, 80.9699, 
    84.04895, 86.31731, 93.66522, 95.5272, 96.60124, 96.82883,
  89.36375, 90.34907, 91.12132, 91.82996, 92.47885, 92.64668, 92.58742, 
    92.35148, 85.8754, 83.96995, 79.57323, 81.56728, 82.41041, 87.29627, 
    88.48795, 82.07735, 82.6252, 91.55006, 89.91431, 91.60603,
  89.04642, 88.77974, 88.9644, 89.50189, 90.48761, 91.16055, 91.46013, 
    91.63289, 89.45311, 89.06082, 88.7837, 88.71642, 88.80796, 89.02697, 
    89.44395, 90.18876, 90.64693, 90.83304, 90.83619, 92.82255,
  91.381, 91.32777, 91.81437, 92.22284, 91.91559, 91.11581, 90.84014, 
    91.22728, 91.88726, 92.61813, 94.01647, 95.52488, 96.17719, 95.62572, 
    94.60149, 93.52795, 92.30692, 91.31403, 90.66068, 90.29609,
  87.94328, 86.93435, 86.53931, 87.45795, 88.3271, 88.51883, 88.52135, 
    89.36317, 90.22198, 91.21557, 92.44796, 93.80112, 94.18541, 93.87446, 
    92.79964, 90.77025, 88.91978, 88.0657, 87.74664, 87.77767,
  87.57671, 86.72248, 85.99305, 86.30566, 87.51836, 88.07648, 87.90142, 
    88.04276, 88.3549, 89.152, 89.43331, 89.50089, 89.58836, 89.9478, 
    90.52554, 90.55193, 89.674, 88.94888, 88.48161, 88.77338,
  91.09366, 90.69493, 89.94524, 89.6131, 89.58879, 88.28461, 85.68106, 
    84.01744, 83.02459, 81.7316, 80.66682, 80.85049, 82.74431, 85.25579, 
    87.15401, 88.78616, 89.61045, 90.03527, 90.19332, 89.97337,
  88.42769, 86.96095, 85.40747, 84.02532, 82.49207, 80.78076, 79.58668, 
    79.1415, 78.64349, 77.87067, 77.23355, 78.19286, 80.47894, 83.30258, 
    85.6786, 87.59331, 87.53833, 87.30034, 87.62063, 88.39135,
  87.44272, 85.1329, 81.59795, 78.95118, 76.53951, 75.15326, 75.37733, 
    76.57459, 77.5612, 78.45411, 79.40772, 81.47527, 84.16791, 85.94182, 
    86.68401, 87.17461, 86.91272, 86.18091, 86.56663, 88.41714,
  83.80001, 81.50262, 76.5315, 73.17826, 72.11286, 73.23222, 75.6178, 
    78.08836, 80.29535, 82.57722, 84.4914, 85.98397, 87.19958, 88.11321, 
    88.24139, 88.11656, 87.58872, 86.67764, 86.82661, 87.35455,
  78.91243, 75.90419, 71.61028, 70.74944, 73.03324, 75.71056, 78.06278, 
    79.94772, 81.68781, 83.4613, 84.88354, 86.16106, 86.99618, 87.57203, 
    87.3634, 86.8417, 85.2104, 83.27094, 81.67094, 80.70864,
  76.79228, 74.66872, 75.24469, 76.88284, 78.40177, 79.45932, 79.43517, 
    76.8298, 74.43923, 74.7774, 76.65799, 79.22164, 81.23644, 81.92094, 
    81.50611, 80.20809, 77.37048, 74.01122, 72.21947, 72.06706,
  76.90186, 78.04296, 78.80404, 78.43445, 77.97784, 75.99397, 70.35272, 
    64.55618, 61.0882, 60.61414, 61.11452, 62.9796, 65.80894, 67.90656, 
    69.76695, 70.35622, 70.04077, 69.70454, 70.13286, 71.1795,
  72.5605, 72.56421, 71.73916, 71.33321, 70.7872, 67.82381, 63.55244, 
    58.4271, 58.62081, 59.94578, 60.73337, 61.85211, 65.73692, 68.172, 
    70.06444, 71.37035, 72.4763, 73.47938, 74.14798, 74.23606,
  92.63737, 92.85606, 92.9079, 93.1693, 93.47414, 93.76683, 93.96848, 
    94.14044, 92.79372, 92.95631, 93.09241, 93.21959, 93.40902, 93.65611, 
    93.78867, 93.81246, 93.02335, 93.12505, 93.25354, 93.10682,
  88.80007, 89.65867, 90.71027, 91.53937, 92.31812, 92.86364, 93.72016, 
    94.43623, 90.77859, 91.4222, 91.98414, 92.27451, 93.03027, 93.40741, 
    93.73303, 93.93841, 91.878, 92.22124, 92.7692, 93.02833,
  85.83212, 87.0879, 88.58112, 90.113, 91.58788, 93.06786, 94.09399, 
    95.10172, 90.94733, 91.78579, 92.2421, 92.40405, 93.47308, 93.77422, 
    94.05655, 94.40392, 91.74497, 92.03923, 92.37429, 92.96049,
  84.81995, 86.21139, 87.36311, 88.5503, 89.65405, 90.58888, 91.64592, 
    92.34897, 89.65915, 90.5115, 91.19485, 91.21816, 91.35768, 91.11637, 
    90.9898, 90.54339, 90.9138, 90.64444, 90.85739, 91.52412,
  83.27023, 85.37543, 87.39245, 89.23051, 90.51286, 91.2197, 91.42264, 
    91.61197, 90.09808, 90.79515, 91.31907, 91.63425, 92.41918, 92.75471, 
    92.67303, 92.64501, 96.92473, 96.84091, 96.34097, 95.686,
  83.35003, 85.97333, 88.1311, 89.62875, 90.57969, 91.19055, 91.32352, 
    91.18848, 87.0349, 87.38918, 88.08676, 89.30901, 90.32298, 91.67606, 
    92.84492, 93.77845, 99.16073, 99.08418, 98.82355, 98.14483,
  89.42117, 86.72526, 85.86785, 86.21218, 86.21551, 86.05222, 86.09634, 
    86.12428, 78.45171, 77.49425, 75.9807, 77.19411, 78.43771, 83.69009, 
    84.33678, 86.17783, 93.67474, 95.59322, 96.65358, 96.9901,
  90.90075, 91.65498, 91.96671, 91.76736, 91.40203, 90.90317, 90.73294, 
    90.12032, 82.37771, 80.06041, 77.28586, 82.49397, 84.08812, 88.64902, 
    79.26662, 76.85034, 76.09283, 92.20461, 92.2989, 93.83093,
  84.8178, 84.50648, 83.60157, 82.35516, 82.25301, 83.22388, 84.10383, 
    83.82995, 80.65698, 80.46426, 81.27192, 82.65815, 84.03626, 84.21373, 
    83.66341, 85.1741, 87.06818, 87.55947, 91.04335, 93.92097,
  81.5846, 81.6426, 82.06268, 79.95638, 77.01954, 75.96516, 75.46899, 
    75.22203, 75.25456, 75.26871, 75.88503, 76.80723, 77.1992, 76.99915, 
    76.4236, 77.07925, 78.35049, 80.68089, 83.39386, 84.84145,
  79.73616, 79.85199, 80.0072, 79.01186, 78.30771, 77.88738, 77.04289, 
    76.2594, 76.53242, 76.85332, 77.59027, 78.41629, 78.02657, 77.03754, 
    76.29731, 76.01929, 76.13636, 77.1072, 78.18671, 79.04147,
  81.3091, 81.37781, 81.16022, 80.67202, 81.09629, 81.85295, 81.44175, 
    80.8069, 80.85204, 81.00898, 80.91855, 81.36843, 81.37039, 80.584, 
    79.13656, 78.9432, 79.5088, 80.02362, 80.20393, 80.9613,
  85.39495, 85.56586, 85.30777, 84.36082, 83.7065, 83.12881, 81.62785, 
    80.93952, 80.52901, 80.38799, 79.73956, 79.97036, 81.57773, 83.60891, 
    84.51754, 85.1347, 84.79665, 84.13165, 83.63648, 83.2167,
  84.92719, 84.27892, 82.7468, 81.06195, 78.44231, 76.87525, 76.91174, 
    77.50268, 78.49165, 79.25893, 79.35128, 80.35293, 82.72083, 85.23074, 
    87.40435, 88.25256, 87.46571, 87.26653, 87.3974, 86.91795,
  84.28381, 82.47392, 79.46979, 77.2003, 75.54485, 74.85, 75.10972, 76.3822, 
    78.34506, 80.06726, 81.39232, 83.38303, 85.96349, 88.21956, 89.08762, 
    89.0355, 88.6983, 88.7306, 89.33891, 90.13624,
  82.33965, 80.25403, 75.27761, 72.41087, 72.29897, 73.425, 75.10864, 
    77.60098, 80.41755, 82.33817, 83.97502, 85.62189, 87.56422, 89.13595, 
    89.05711, 88.54465, 87.86732, 87.44813, 88.15701, 88.62633,
  78.12691, 75.96215, 72.96832, 71.96037, 73.13195, 74.70911, 76.39874, 
    77.83069, 79.43853, 81.15201, 82.64734, 83.75937, 84.66048, 85.46927, 
    85.37489, 84.61079, 82.992, 81.74709, 81.16718, 80.54422,
  74.62702, 73.57899, 73.97563, 75.37119, 77.25686, 78.3002, 78.20376, 
    76.1405, 73.38818, 73.03576, 74.45078, 76.77982, 78.84028, 79.51389, 
    79.48599, 78.45872, 75.13653, 71.70178, 70.25199, 70.72385,
  72.24899, 73.71836, 75.0655, 75.48645, 76.07313, 75.35955, 72.02425, 
    66.39941, 61.21125, 59.39012, 60.81732, 63.06049, 65.86478, 67.96339, 
    68.9578, 68.86578, 67.83147, 67.38908, 68.43168, 69.92563,
  68.46617, 69.2587, 68.79629, 69.03622, 69.83079, 68.31286, 65.85081, 
    61.7156, 60.24652, 59.74588, 62.38418, 64.07027, 67.29463, 69.35155, 
    69.86797, 70.33462, 70.67255, 71.08336, 71.69938, 71.6804,
  89.36323, 89.58965, 89.93466, 90.11516, 90.33382, 90.6096, 90.94618, 
    91.226, 89.71793, 89.88908, 90.08227, 90.36639, 90.51334, 90.82721, 
    91.15472, 91.77075, 91.16086, 91.08852, 91.47682, 91.80979,
  85.55634, 86.51617, 87.45711, 88.3218, 89.28326, 90.1478, 91.10569, 
    92.0163, 88.58524, 89.42967, 90.14968, 90.79809, 91.53135, 92.30772, 
    93.14343, 93.91769, 92.05259, 92.68748, 93.50358, 94.16422,
  86.19411, 87.46588, 88.76097, 89.92612, 91.12273, 92.31626, 93.4525, 
    94.40907, 90.07473, 91.16891, 92.45821, 93.68399, 94.58664, 95.5007, 
    96.23571, 97.03107, 95.63757, 96.04101, 96.46251, 96.91166,
  87.19146, 88.59389, 90.22549, 91.77813, 92.79789, 93.70517, 94.39866, 
    94.88293, 92.30849, 93.00256, 94.01151, 94.94733, 95.77652, 96.64886, 
    97.41837, 97.79739, 98.50916, 98.54092, 98.38778, 98.14349,
  86.47557, 88.04025, 88.4994, 89.02061, 90.7451, 91.97108, 93.0566, 
    93.93545, 93.20985, 93.6829, 94.40501, 95.21008, 95.69959, 96.30609, 
    96.90161, 97.13321, 99.33077, 99.12022, 98.54219, 97.81819,
  83.4453, 85.55761, 87.08728, 88.2672, 89.22458, 89.75143, 89.62032, 
    89.93008, 85.91712, 86.72665, 87.54719, 88.6775, 89.82661, 91.04811, 
    92.5334, 93.69405, 98.63773, 98.63972, 98.35879, 97.7314,
  91.09675, 88.9903, 87.60851, 87.23551, 87.12933, 87.84913, 88.51283, 
    88.61292, 80.82629, 79.82373, 78.51551, 76.55662, 78.6287, 87.01571, 
    90.22678, 84.90505, 92.22346, 95.07462, 96.56784, 96.75105,
  75.52678, 74.82759, 73.47547, 72.00417, 72.3222, 73.33171, 73.32531, 
    72.44235, 65.27482, 63.35582, 63.43764, 71.12511, 70.80512, 76.0398, 
    71.5564, 73.80165, 84.23235, 90.31237, 87.16445, 89.00074,
  73.89975, 74.14558, 74.7594, 75.61689, 77.42399, 79.75613, 81.77088, 
    82.81993, 80.73122, 80.51241, 79.68671, 78.0448, 75.93897, 72.93349, 
    70.72813, 71.80161, 72.41516, 71.1395, 77.09783, 79.19968,
  76.16766, 76.32806, 76.97137, 77.55979, 77.69455, 78.72591, 80.50827, 
    82.47748, 83.68138, 84.53767, 85.27789, 85.25313, 83.76477, 81.53177, 
    78.58308, 76.37331, 75.83833, 77.06728, 78.59396, 79.5114,
  78.98853, 78.42474, 78.65466, 79.12992, 80.06923, 80.96443, 81.45782, 
    82.62399, 83.40668, 84.58566, 85.99611, 87.27935, 87.05808, 85.47914, 
    83.75832, 82.16619, 81.84159, 82.47732, 83.68394, 84.83515,
  84.10291, 83.09241, 82.34934, 82.2439, 82.45776, 82.29217, 81.90427, 
    82.70459, 84.07742, 85.55709, 86.44476, 87.42266, 88.39068, 88.3626, 
    87.70622, 87.50019, 88.59536, 89.52209, 89.78574, 89.81654,
  87.24152, 86.99991, 86.82542, 86.2019, 84.81346, 83.16975, 81.55824, 
    81.52905, 82.38771, 83.10915, 83.64405, 84.4861, 86.31034, 88.72421, 
    90.88197, 92.58135, 93.78683, 94.32088, 94.15279, 93.12746,
  86.00883, 85.1715, 84.23861, 83.4494, 82.26853, 81.26782, 80.47736, 
    80.33094, 81.04366, 81.90851, 82.95253, 84.60819, 86.91918, 89.49025, 
    92.1236, 93.98371, 94.13464, 93.97292, 94.18387, 93.90679,
  86.9512, 84.90179, 82.49248, 80.71213, 78.93139, 78.08192, 78.27573, 
    79.07906, 80.61844, 82.38902, 84.12449, 86.08372, 88.17793, 90.04402, 
    91.76836, 92.61362, 92.58506, 92.45403, 92.92478, 93.5329,
  84.63981, 82.46618, 78.77744, 76.96116, 76.64273, 77.84743, 79.92317, 
    81.67298, 83.21587, 84.6665, 85.96346, 87.36695, 88.71542, 89.93964, 
    90.04819, 89.85242, 90.24272, 90.6256, 91.27043, 91.12238,
  79.65468, 78.11831, 77.38485, 78.51028, 79.43709, 80.79626, 81.64131, 
    82.01329, 82.82668, 83.55342, 84.24686, 84.97982, 85.77937, 86.13979, 
    86.16843, 86.17906, 86.01617, 85.7366, 85.57327, 85.9876,
  78.82792, 78.88149, 79.67372, 80.52344, 80.61268, 79.78967, 78.02666, 
    75.83865, 74.40656, 74.74137, 75.72167, 77.16711, 79.23126, 81.15778, 
    82.19939, 82.65479, 81.97025, 80.64296, 80.95997, 82.39488,
  78.23505, 77.60584, 76.6049, 75.15005, 74.37511, 72.65833, 69.80402, 
    66.73027, 64.19173, 63.5056, 63.2512, 64.64748, 67.93256, 71.39038, 
    74.67421, 76.40465, 77.41135, 77.46899, 78.64718, 79.49009,
  72.23376, 71.0588, 69.34719, 69.03336, 70.80698, 70.91716, 70.49986, 
    68.75531, 68.60476, 69.36029, 67.99298, 67.64799, 70.72482, 73.24512, 
    75.39919, 77.56806, 78.97816, 79.27144, 79.04144, 77.12852,
  91.23755, 91.65125, 92.12211, 92.6165, 93.1147, 93.42018, 93.94121, 
    94.32806, 93.0918, 93.54514, 93.83637, 94.20033, 94.46982, 94.72564, 
    95.16801, 95.25451, 94.38379, 94.58986, 94.89684, 95.06989,
  85.86654, 87.19549, 88.51644, 89.79427, 90.97515, 91.90726, 92.76971, 
    93.53024, 90.15945, 91.25708, 92.42744, 93.58237, 94.45453, 95.08404, 
    95.7157, 95.91708, 94.31877, 94.84076, 95.28856, 95.70432,
  85.945, 87.67599, 89.33908, 90.58085, 91.86753, 93.16286, 93.91825, 
    94.48253, 90.21141, 91.00108, 91.83501, 93.06914, 94.52168, 95.92642, 
    97.15137, 98.14687, 97.18304, 97.77951, 98.01721, 98.28638,
  84.94824, 86.44317, 87.93915, 89.43398, 90.56267, 91.44783, 92.03454, 
    92.29791, 89.70676, 90.50259, 92.75861, 95.07896, 96.90237, 98.08536, 
    98.93497, 99.1468, 99.52171, 99.54363, 99.39876, 99.21582,
  82.72894, 83.79469, 85.02325, 85.35605, 84.49635, 83.86371, 83.66322, 
    83.53263, 83.47572, 85.54064, 87.71006, 90.15694, 92.68309, 94.75833, 
    95.84998, 96.22226, 98.74629, 98.72772, 98.42733, 97.92953,
  79.75217, 82.13435, 84.16023, 85.2179, 85.71957, 85.84035, 85.88818, 
    85.94701, 82.14114, 82.60937, 83.46783, 84.81229, 86.50163, 87.87977, 
    88.9007, 89.39877, 95.75515, 96.20937, 96.22384, 95.88781,
  90.99618, 90.51688, 90.62746, 90.75703, 91.09086, 91.69654, 92.13428, 
    92.33716, 84.85445, 84.92754, 84.41753, 76.75642, 78.37951, 85.02744, 
    88.37991, 85.01358, 91.31927, 93.55349, 95.03269, 95.30099,
  76.5184, 76.47433, 75.97572, 76.02338, 77.26179, 80.68526, 79.15479, 
    77.79886, 68.91508, 66.70721, 65.5084, 68.92612, 74.13354, 82.85302, 
    86.65831, 88.05072, 90.90915, 89.95197, 86.94922, 85.40303,
  75.87701, 74.58003, 73.05978, 71.67186, 70.80466, 70.37325, 70.07575, 
    69.47612, 66.38763, 65.98209, 65.3, 64.93398, 65.90826, 67.62041, 
    69.44299, 71.71364, 73.89096, 76.65171, 80.5631, 84.0473,
  75.84319, 76.34981, 76.68953, 76.80045, 76.43673, 76.0469, 75.93713, 
    75.60265, 75.20849, 75.00204, 74.44897, 73.87041, 73.66396, 73.60966, 
    73.28785, 73.85635, 75.36977, 76.91047, 78.06101, 77.93257,
  78.03769, 77.26905, 77.36642, 78.40619, 79.19623, 79.42538, 79.56855, 
    79.84435, 80.02773, 79.9418, 79.79518, 79.60674, 79.42854, 79.26006, 
    79.76618, 80.39294, 81.57636, 82.71894, 83.57541, 84.53719,
  82.24799, 80.42308, 79.50498, 79.31488, 79.30357, 78.72606, 78.43129, 
    79.24343, 80.64642, 81.7091, 82.05409, 82.17147, 82.58917, 83.36646, 
    84.0647, 84.1353, 84.45689, 85.11906, 85.1309, 85.33992,
  85.09152, 83.62634, 82.5863, 82.04299, 81.12962, 79.33567, 77.22773, 
    76.25695, 76.19583, 76.7329, 77.29982, 78.01664, 78.93098, 80.54357, 
    82.68613, 84.1842, 85.25536, 85.84605, 86.08891, 85.31341,
  83.54884, 81.8567, 80.11267, 79.10838, 77.9314, 76.44716, 75.22559, 
    74.36304, 73.73615, 73.67086, 73.97129, 74.79317, 76.51524, 78.9828, 
    81.58358, 83.87946, 85.21647, 86.44876, 87.73447, 88.41785,
  83.48231, 81.35819, 78.42453, 76.51283, 74.73693, 73.44465, 73.00938, 
    73.17562, 73.23306, 73.77105, 74.86565, 76.60387, 78.64862, 80.79995, 
    82.2337, 83.48605, 84.55688, 85.55563, 87.15588, 88.76123,
  83.45997, 80.89696, 76.27486, 73.85138, 73.77387, 74.48, 74.97176, 
    76.10352, 77.06294, 78.09113, 79.03375, 79.97018, 80.91047, 81.64262, 
    81.73473, 81.73495, 81.62822, 81.44468, 82.42255, 83.43884,
  82.16373, 79.00035, 76.60954, 76.96187, 78.52971, 79.54368, 79.6962, 
    78.81583, 78.07265, 78.14142, 78.83212, 79.57205, 79.97585, 79.56664, 
    78.35145, 77.34664, 76.16398, 74.55747, 73.70211, 74.03942,
  81.47728, 80.22129, 80.6217, 81.07948, 81.34439, 80.47222, 77.27724, 
    71.77167, 67.60878, 67.52163, 69.30412, 71.41422, 72.40205, 71.5303, 
    70.92034, 70.9315, 69.61764, 67.66959, 67.39905, 68.41116,
  76.93097, 77.00003, 76.45455, 74.80365, 73.69473, 72.0807, 67.98618, 
    63.33226, 60.85281, 60.3437, 60.704, 60.85299, 62.04815, 63.50024, 
    64.62486, 65.08096, 65.63734, 66.43282, 67.74477, 68.55895,
  68.57254, 68.12991, 66.79195, 66.4548, 68.58408, 69.87177, 70.79552, 
    69.11112, 69.0018, 68.29599, 66.7558, 65.39233, 66.98226, 68.57095, 
    68.47585, 68.2534, 68.4782, 69.31599, 70.45207, 70.46724,
  93.33907, 93.68111, 94.00677, 94.19484, 94.54321, 94.96457, 95.19604, 
    95.38432, 94.11292, 94.68447, 94.87923, 94.99619, 95.37181, 95.74664, 
    96.07202, 96.66339, 96.08672, 96.78719, 97.43752, 97.77699,
  86.92452, 87.92088, 88.86559, 89.77613, 90.65554, 91.67281, 92.94258, 
    94.08537, 90.93831, 92.45257, 93.43297, 94.30183, 95.05526, 95.89188, 
    96.44382, 96.89111, 95.85049, 96.35027, 96.78364, 97.67533,
  86.75605, 88.28974, 89.49566, 90.66571, 92.14505, 93.53957, 94.54973, 
    95.91028, 91.78979, 93.02241, 93.87985, 94.66617, 95.36656, 95.98984, 
    96.56336, 96.82375, 96.67851, 97.85739, 98.46918, 99.00564,
  83.25169, 85.69691, 87.78256, 89.45901, 90.5836, 91.81833, 93.4329, 
    94.97913, 94.2412, 95.38906, 96.37039, 97.50417, 98.36926, 99.07334, 
    99.37759, 99.32133, 99.50452, 99.74392, 99.68085, 99.27176,
  77.04681, 79.39981, 80.82032, 81.61044, 81.70638, 82.53448, 83.96849, 
    85.75833, 86.11182, 88.63568, 91.31161, 93.55354, 95.1105, 95.90039, 
    95.92458, 96.02366, 98.33645, 98.43318, 98.38544, 97.9793,
  78.86657, 79.04941, 80.20735, 81.18478, 81.60722, 81.7077, 82.58453, 
    83.08841, 79.94435, 81.17639, 82.44353, 83.80031, 84.91951, 85.80936, 
    86.04352, 86.48412, 93.02023, 93.7144, 94.08289, 93.75498,
  89.81462, 86.49056, 86.89929, 88.03967, 88.95261, 88.89403, 88.01462, 
    87.34591, 80.26913, 81.56844, 83.86753, 75.93755, 78.26119, 85.70664, 
    89.63199, 86.06947, 91.8928, 93.0757, 94.24819, 93.97298,
  88.07516, 86.44093, 84.43246, 83.97398, 84.27536, 85.13602, 85.52676, 
    86.16151, 81.24619, 83.70393, 87.18151, 83.5455, 85.03626, 91.0948, 
    93.3923, 96.31415, 97.30685, 94.89188, 92.30175, 92.2859,
  68.768, 66.4192, 65.03826, 64.34743, 64.60775, 66.11805, 66.34441, 
    65.78966, 63.87374, 63.48436, 62.40854, 63.87227, 69.7599, 75.8205, 
    80.99976, 84.99221, 88.63824, 92.28506, 94.74667, 95.73791,
  76.99828, 76.15809, 75.43842, 74.68504, 74.10041, 73.74654, 73.19926, 
    72.56258, 72.48438, 72.34859, 71.78754, 70.64801, 70.40578, 70.44646, 
    70.45025, 70.93952, 72.40169, 73.43736, 74.43226, 75.33275,
  80.63052, 79.87993, 79.46091, 79.08664, 78.70894, 78.36465, 78.1549, 
    78.04682, 78.53964, 78.84249, 78.95396, 79.09467, 79.4187, 79.77305, 
    80.17607, 80.68182, 81.24084, 80.86668, 80.38146, 79.90677,
  83.61308, 83.29057, 83.22675, 83.39452, 83.37061, 82.80448, 82.09825, 
    82.5153, 83.64931, 83.45671, 82.52151, 82.04947, 82.79562, 83.80991, 
    84.76179, 85.27483, 86.29817, 86.68304, 86.34251, 85.51234,
  87.1746, 87.09988, 87.04337, 86.9765, 86.46247, 84.55501, 82.01046, 
    80.54957, 79.90945, 79.27916, 79.03314, 79.88095, 82.01077, 84.34393, 
    86.59843, 88.65417, 90.28941, 90.61062, 90.19366, 88.91532,
  83.92834, 82.39164, 80.79478, 79.34028, 77.71048, 76.60547, 76.07832, 
    76.10722, 77.08892, 78.41495, 79.86176, 81.64085, 84.22253, 87.29054, 
    89.77778, 91.50121, 92.22177, 92.15589, 91.97823, 91.73212,
  81.28149, 78.29086, 74.58802, 71.57955, 68.99265, 68.30982, 69.41199, 
    71.40435, 74.46632, 77.39032, 80.23703, 83.36365, 86.28221, 88.58372, 
    89.92451, 90.4226, 90.41959, 89.79176, 90.07088, 91.07803,
  76.19399, 73.0272, 67.1848, 63.95276, 63.91945, 65.95623, 68.35077, 
    71.25965, 75.35279, 79.46268, 83.0768, 85.32672, 86.95812, 88.29709, 
    88.521, 87.98049, 87.2551, 86.39385, 87.00076, 87.83495,
  67.28919, 63.57757, 61.72634, 63.40101, 66.16788, 69.11356, 71.46201, 
    73.65742, 76.31405, 79.28497, 81.67857, 83.73277, 85.70283, 86.83546, 
    86.63546, 85.14453, 83.17761, 81.52481, 81.21373, 81.32195,
  63.78304, 63.86884, 66.18721, 68.73483, 70.24429, 70.32754, 68.86571, 
    64.5416, 61.45775, 61.99194, 65.4419, 71.21131, 77.41018, 80.99164, 
    81.77641, 80.78315, 78.41146, 75.89075, 74.75375, 74.00346,
  67.47063, 69.56741, 70.62238, 69.24794, 67.13795, 64.09286, 58.86689, 
    54.41287, 53.59605, 53.83799, 54.96211, 58.55197, 63.04151, 67.41283, 
    71.44672, 72.99784, 73.3242, 72.63551, 72.14408, 71.96929,
  64.92885, 65.47015, 64.41721, 62.69117, 62.02641, 60.79371, 61.4697, 
    61.26355, 61.68913, 62.62842, 61.34033, 62.30093, 65.61166, 69.84261, 
    73.30482, 75.01622, 75.39145, 74.76627, 74.12801, 72.64287,
  90.052, 90.56416, 91.06026, 91.61353, 92.02836, 92.40627, 92.78955, 
    93.14735, 92.00945, 92.31061, 92.58345, 92.99615, 93.28033, 93.57104, 
    93.76012, 94.04841, 93.38367, 93.34415, 93.54231, 93.55079,
  86.97238, 88.54171, 89.96096, 91.40443, 92.70685, 93.8036, 94.61906, 
    95.44979, 92.20555, 93.05804, 93.86304, 94.53702, 95.27808, 96.12707, 
    96.84732, 97.59583, 96.11971, 96.59029, 96.77213, 96.93997,
  83.69521, 85.69416, 87.72955, 89.86126, 91.78108, 93.55563, 94.96161, 
    96.27407, 92.37347, 92.97688, 94.23998, 95.34776, 96.64389, 97.86816, 
    98.69823, 98.65619, 98.25706, 98.31248, 98.19617, 98.34538,
  85.3348, 88.12923, 90.63098, 92.6326, 94.54549, 95.85041, 96.54823, 
    96.91792, 94.70312, 95.78383, 97.35541, 98.2319, 98.6749, 98.6244, 
    98.79445, 98.95319, 99.05836, 99.12052, 99.00632, 98.56697,
  83.29901, 86.50014, 89.08883, 90.26991, 91.4087, 92.44244, 93.0614, 
    93.98579, 93.95943, 94.90604, 94.62608, 95.21797, 96.24723, 96.51029, 
    96.82793, 97.53316, 98.98804, 99.10126, 99.33981, 98.51507,
  80.15831, 81.2654, 82.86002, 83.88515, 84.45975, 85.10019, 85.71247, 
    86.57873, 83.17428, 83.1588, 82.90812, 84.02054, 85.30446, 86.7434, 
    88.08796, 89.70208, 94.65679, 95.82561, 96.88232, 97.46455,
  94.19733, 89.60251, 89.5726, 89.84374, 89.93987, 89.71503, 89.03501, 
    88.48397, 80.58302, 81.29348, 83.80947, 74.75541, 77.00272, 84.53638, 
    88.29975, 83.94041, 89.89257, 91.27498, 92.59669, 93.50683,
  95.99648, 95.29808, 94.72274, 94.32397, 94.2173, 95.0213, 95.30936, 
    94.88113, 90.47065, 91.73029, 93.76001, 89.14172, 89.98575, 92.76893, 
    95.10273, 96.45982, 97.05594, 95.68123, 93.08547, 93.06852,
  95.45928, 94.27051, 93.32242, 93.42924, 94.47848, 95.50489, 95.63498, 
    95.57008, 94.26073, 94.28156, 94.46203, 94.80473, 94.13033, 93.62237, 
    92.40672, 91.6082, 93.81405, 96.52575, 97.41669, 95.68252,
  74.88612, 74.72481, 73.48712, 73.22332, 74.71289, 77.64471, 80.07373, 
    80.58073, 79.75966, 77.14314, 75.04176, 74.51174, 75.42038, 75.85256, 
    74.85125, 74.99477, 76.57569, 80.46826, 85.81409, 89.46384,
  61.50371, 61.66653, 61.33796, 61.14944, 61.36743, 62.76193, 64.95052, 
    67.27765, 68.59892, 68.37923, 68.28425, 68.65185, 69.10056, 69.37196, 
    69.58539, 69.97968, 70.91395, 71.88103, 73.13647, 74.30247,
  62.64985, 62.82164, 63.11253, 63.82331, 64.50051, 64.7811, 65.62944, 
    68.08525, 70.55974, 71.76437, 72.47199, 73.25343, 74.35408, 75.58877, 
    76.28449, 76.54095, 77.25966, 77.89943, 77.66528, 76.69373,
  68.42458, 68.03608, 68.07262, 68.34755, 68.25082, 67.29825, 66.64023, 
    67.46102, 69.21513, 70.60555, 71.20954, 71.8418, 72.99478, 75.0357, 
    77.38499, 79.24842, 80.64129, 80.53452, 79.31378, 77.52521,
  73.5392, 71.8535, 70.17406, 68.85921, 67.3191, 66.04506, 66.08419, 
    67.38422, 69.09852, 70.42355, 71.14944, 71.77791, 72.45866, 74.84406, 
    78.40359, 80.75378, 81.38392, 81.22253, 80.92377, 80.02032,
  75.74944, 73.61049, 70.80848, 68.10119, 65.24911, 63.63064, 64.17072, 
    66.13307, 68.83073, 71.33078, 73.34187, 75.12338, 76.89085, 79.08035, 
    81.49112, 83.05952, 83.234, 82.35979, 81.64119, 81.55163,
  76.16044, 74.06783, 69.02173, 64.7591, 63.25753, 64.27224, 66.88486, 
    69.90324, 73.59926, 76.82942, 79.37724, 81.31844, 82.94897, 84.3194, 
    84.64285, 84.04813, 82.31074, 80.22932, 79.72982, 79.93727,
  73.26598, 70.29649, 67.73515, 68.57722, 70.53045, 73.11925, 75.95997, 
    78.4422, 80.52903, 82.38853, 83.90744, 84.86803, 85.11133, 84.93281, 
    83.8916, 82.15507, 79.13519, 75.83009, 73.65845, 73.32755,
  69.70096, 71.06816, 74.47994, 77.35672, 78.85219, 79.25265, 77.58596, 
    72.79974, 68.88995, 68.72219, 71.33065, 75.258, 78.61165, 79.84354, 
    79.27828, 77.7182, 74.01077, 69.90995, 67.92748, 68.45056,
  68.07788, 71.54037, 74.33728, 74.35297, 73.76237, 71.1835, 65.71567, 
    61.07678, 59.79924, 58.96383, 59.46315, 61.9069, 65.37065, 67.78869, 
    68.26717, 67.79836, 67.37128, 67.8217, 69.30281, 71.17813,
  63.24943, 65.18267, 66.30532, 66.63465, 66.89183, 66.24466, 65.48817, 
    65.06051, 65.86863, 64.78381, 61.1033, 61.61998, 66.21956, 69.99608, 
    70.43285, 70.26716, 70.88605, 72.34962, 74.03788, 74.93484,
  93.15509, 93.45945, 94.04833, 94.38045, 94.81377, 95.31415, 95.61769, 
    95.95625, 95.01917, 95.78452, 96.06263, 96.6142, 96.81416, 97.21481, 
    97.13115, 97.59377, 97.02632, 97.13256, 97.14542, 97.09566,
  86.51275, 88.03004, 89.5089, 90.96017, 92.28883, 93.37366, 94.04926, 
    94.80756, 91.31112, 91.76744, 92.12809, 93.89271, 94.69435, 95.58411, 
    96.18114, 96.63713, 95.83125, 96.66775, 97.22347, 97.85841,
  89.48326, 91.42107, 93.00645, 94.30444, 95.20441, 95.60303, 95.65044, 
    96.19363, 91.48202, 91.96961, 93.37182, 94.83141, 96.57045, 97.6682, 
    98.46512, 98.89157, 98.68521, 99.33546, 99.74779, 99.92838,
  89.5395, 91.48708, 93.05704, 94.13654, 95.44892, 96.59918, 97.83035, 
    98.58327, 97.19698, 96.97444, 97.30101, 97.73955, 98.83945, 99.41248, 
    99.74586, 99.83145, 99.84642, 99.85196, 99.87671, 99.83685,
  87.27375, 90.52389, 92.75864, 93.99734, 94.54557, 93.33199, 92.68354, 
    93.00479, 92.43794, 91.51383, 91.48959, 92.06098, 93.18015, 94.70052, 
    96.19336, 97.49991, 99.19305, 99.34774, 99.3252, 99.21825,
  82.66785, 84.74672, 86.25427, 87.04249, 86.70742, 86.37138, 87.06366, 
    88.00148, 83.93501, 84.1254, 84.60705, 85.52911, 86.73483, 88.11993, 
    89.62698, 91.09261, 96.99282, 97.67976, 98.16284, 98.68069,
  96.70408, 91.83814, 90.76633, 90.64675, 90.14999, 89.38017, 87.92052, 
    87.34032, 79.59825, 81.00829, 83.62798, 76.48495, 77.87923, 83.67704, 
    87.85438, 84.02428, 90.38895, 92.49608, 93.78462, 94.52805,
  97.54564, 97.46192, 97.28527, 97.29749, 96.75423, 96.59406, 95.96805, 
    95.27711, 90.84038, 91.67432, 92.93423, 87.3921, 88.40701, 93.25792, 
    96.3941, 95.32647, 95.901, 93.04374, 89.43114, 89.83405,
  97.32135, 96.98945, 96.65236, 97.48735, 98.56217, 98.7136, 98.33202, 
    97.73898, 95.36314, 95.22313, 95.6, 96.47247, 96.75701, 97.11259, 
    96.88796, 97.23771, 98.44875, 98.85201, 99.07498, 98.54417,
  96.68538, 96.10732, 96.42233, 97.00667, 97.47537, 97.10028, 96.56441, 
    95.8863, 94.52483, 94.59132, 95.37372, 96.30593, 96.6589, 96.09449, 
    94.59914, 94.26075, 94.35641, 94.67485, 96.01647, 96.82957,
  94.9968, 95.24927, 94.75831, 95.14489, 93.59846, 89.03542, 85.47945, 
    84.82906, 84.66155, 84.4733, 83.76083, 83.54044, 84.14412, 84.49907, 
    83.05495, 80.00546, 76.82607, 72.65164, 68.62318, 67.71835,
  77.70366, 77.43629, 75.90578, 75.52489, 74.08781, 69.88177, 66.46507, 
    66.40284, 67.40018, 68.02547, 68.41896, 68.80045, 69.55831, 70.76044, 
    71.97243, 72.29853, 72.83424, 72.99352, 71.86417, 69.57412,
  77.91448, 77.42785, 77.04996, 76.58544, 75.4646, 73.41133, 71.3075, 
    70.6416, 71.14767, 71.71026, 71.52028, 70.93884, 70.68832, 71.48521, 
    73.26675, 74.93056, 76.47382, 77.44771, 77.28885, 76.3615,
  80.89172, 79.37794, 77.61389, 75.95087, 74.0694, 72.6936, 72.23232, 
    72.51211, 72.9338, 72.855, 72.27521, 71.99015, 72.25356, 73.68248, 
    76.66882, 78.99599, 79.7257, 80.29941, 81.30636, 82.20962,
  81.16671, 78.58562, 74.83076, 71.95668, 69.4791, 68.10172, 68.56696, 
    69.98441, 71.04376, 71.91601, 72.82556, 74.29292, 75.9398, 77.51922, 
    79.45837, 80.92579, 81.6537, 81.99884, 83.00166, 84.72372,
  79.8616, 77.27617, 70.94536, 66.25591, 64.52091, 65.21459, 67.74541, 
    70.82401, 73.59471, 76.27961, 78.66975, 80.31213, 81.53217, 82.71806, 
    83.45065, 83.71896, 83.36841, 82.50745, 83.07975, 84.42816,
  75.51318, 70.81417, 66.18764, 65.93736, 67.66396, 70.38816, 74.07508, 
    77.43066, 79.82453, 81.69041, 82.96809, 83.77124, 84.09564, 84.37923, 
    84.51466, 84.11797, 82.31886, 80.06226, 78.45016, 77.53828,
  69.87688, 69.26967, 71.21701, 73.7653, 75.88224, 77.64854, 76.9507, 
    72.65964, 69.05386, 68.53112, 70.13106, 73.3382, 76.61799, 78.31525, 
    78.63985, 77.38747, 73.61626, 69.03445, 66.83358, 66.12276,
  71.66061, 73.79192, 75.33561, 75.08233, 74.60169, 71.80068, 65.87996, 
    60.76789, 59.19752, 56.98579, 55.81915, 56.2434, 58.09644, 60.04312, 
    60.98159, 60.88643, 60.54443, 60.62257, 61.63421, 63.16565,
  69.98058, 70.23722, 69.72493, 69.58389, 69.42001, 67.44389, 65.76846, 
    68.07301, 68.23441, 64.95541, 58.43159, 56.25373, 58.79282, 61.30151, 
    61.79278, 62.1861, 63.50285, 65.23103, 67.32514, 69.36961,
  92.69642, 93.02699, 93.23515, 93.47101, 93.97298, 94.55976, 94.94784, 
    95.34948, 93.99782, 94.55984, 94.89692, 95.22736, 95.5579, 95.93532, 
    96.14516, 96.30161, 95.67522, 95.86275, 96.0777, 96.19814,
  88.05411, 89.15829, 90.29722, 91.48946, 92.69419, 93.91643, 94.89613, 
    95.85819, 92.90344, 93.19262, 93.62348, 94.18838, 94.80737, 95.63248, 
    96.12798, 96.41041, 95.0844, 95.52985, 95.93182, 96.40731,
  88.85448, 90.64867, 92.04226, 93.17001, 94.13261, 94.83712, 95.32655, 
    95.81812, 90.76302, 91.399, 92.65466, 94.76667, 96.24706, 97.19792, 
    97.68725, 98.09511, 97.68633, 98.40942, 98.86411, 99.17112,
  89.58559, 90.9627, 92.16225, 93.09254, 94.33893, 95.52541, 96.36195, 
    96.95253, 95.45553, 96.18459, 96.63586, 97.09889, 97.56619, 98.16265, 
    99.08279, 99.42054, 99.73486, 99.82499, 99.82818, 99.5109,
  87.47525, 89.01035, 90.29819, 91.33223, 92.47147, 93.80567, 94.50476, 
    94.7698, 93.50892, 94.04343, 93.97147, 93.86729, 93.52602, 94.09066, 
    94.76733, 95.13254, 96.93384, 97.60445, 97.88661, 98.47488,
  83.79855, 85.81705, 87.27676, 88.45628, 89.20399, 90.2841, 90.99754, 
    91.03114, 86.12614, 86.11866, 86.38046, 86.92978, 87.45721, 87.2361, 
    87.07339, 87.53088, 92.90876, 95.00202, 96.2339, 96.65466,
  96.35281, 93.94097, 94.37543, 94.58118, 93.73057, 93.8135, 93.38744, 
    91.9817, 83.07423, 81.91545, 81.42699, 75.29072, 76.59237, 83.93899, 
    83.82659, 79.36124, 87.15455, 90.04865, 91.37505, 91.8819,
  98.97772, 99.2271, 99.23423, 98.57838, 98.32172, 99.35439, 99.07899, 
    98.85641, 94.02381, 93.33766, 93.33151, 92.28548, 91.72341, 93.0721, 
    94.17262, 88.46051, 90.59057, 91.25916, 83.54655, 84.54344,
  98.24734, 98.35376, 98.22073, 97.51282, 96.78201, 96.50089, 97.2163, 
    97.24603, 96.06899, 96.30357, 95.99774, 95.86075, 96.01965, 96.08869, 
    96.58699, 96.35844, 95.99557, 96.62055, 96.62363, 96.88275,
  97.01999, 96.72365, 96.75586, 96.83725, 96.32251, 95.24567, 94.26084, 
    94.57573, 95.72977, 96.29572, 96.47234, 96.35031, 96.17508, 96.43655, 
    97.16208, 97.06121, 96.21195, 95.80374, 96.01478, 96.78935,
  95.85925, 95.54188, 95.26398, 94.81905, 94.54916, 94.62911, 93.40559, 
    92.79895, 92.72781, 92.73705, 92.66735, 93.17702, 93.81258, 94.3511, 
    95.26188, 95.33497, 94.7392, 93.98393, 90.47628, 85.7281,
  92.30613, 90.66506, 89.89359, 88.62733, 88.19055, 83.27531, 77.05272, 
    74.8377, 74.24136, 73.78212, 72.67384, 71.98675, 72.63828, 74.47156, 
    75.91018, 76.50541, 78.47594, 79.16582, 71.47587, 63.09346,
  78.38456, 77.86618, 77.97152, 78.71314, 78.8115, 77.8559, 76.63132, 
    76.12202, 76.31337, 75.92548, 74.81804, 73.32766, 71.94121, 71.22514, 
    71.34202, 71.9015, 71.36993, 70.39249, 68.43142, 65.95586,
  81.38535, 81.42634, 81.13518, 80.54855, 79.44202, 78.2373, 77.47458, 
    77.23296, 77.17494, 77.81328, 77.87826, 77.6092, 77.01514, 76.49104, 
    76.65121, 77.07774, 75.93315, 75.09224, 74.68379, 74.24256,
  81.43556, 80.90685, 78.91106, 77.05393, 75.50421, 74.30585, 73.51998, 
    73.14249, 73.10081, 74.14355, 75.33359, 76.85178, 77.91405, 78.20579, 
    78.39954, 78.92513, 78.36527, 78.17402, 78.60346, 79.32494,
  77.84129, 77.59418, 74.34034, 71.19804, 69.55954, 69.29985, 69.41768, 
    70.10696, 71.3988, 73.24528, 75.48204, 77.46036, 78.87718, 80.18053, 
    80.53161, 80.30567, 78.91698, 77.59673, 77.58672, 77.82059,
  70.72034, 68.46133, 64.38342, 64.61651, 67.0878, 69.19292, 71.06405, 
    73.0524, 74.48219, 75.73045, 76.97406, 78.13201, 79.38383, 80.27711, 
    79.58229, 77.96455, 74.94609, 72.22891, 70.61666, 69.88404,
  61.98864, 64.24064, 68.62841, 72.57996, 75.71281, 77.65537, 76.96146, 
    72.07191, 67.57525, 65.99017, 66.29475, 68.04552, 70.46638, 71.80997, 
    71.85954, 70.6573, 66.79012, 62.71004, 61.12037, 61.65081,
  67.51369, 72.44603, 75.56437, 76.98877, 77.16618, 74.03388, 67.77511, 
    62.87537, 60.90215, 58.32723, 57.31681, 57.90615, 59.06445, 59.38869, 
    59.13268, 58.31083, 57.20226, 57.32901, 58.78182, 60.60358,
  69.30038, 70.21964, 70.08711, 70.70155, 69.60519, 66.32713, 64.89326, 
    68.93518, 69.80039, 67.26402, 60.45775, 58.27094, 61.55651, 62.62687, 
    60.34216, 59.11612, 59.99855, 61.76248, 63.38121, 64.90251,
  89.38627, 89.92767, 90.19828, 90.61964, 91.29128, 91.72019, 92.42922, 
    92.71449, 91.58955, 91.97433, 92.36914, 92.7503, 93.26569, 93.70335, 
    94.08855, 94.43033, 93.82826, 94.15947, 94.42857, 94.86898,
  83.68914, 85.29691, 86.82805, 88.44012, 90.04511, 91.5343, 92.76714, 
    93.82818, 90.36461, 90.87021, 91.59927, 91.63394, 92.12609, 92.96471, 
    93.7253, 94.34848, 93.08196, 93.90517, 94.80445, 95.4052,
  84.94196, 86.68272, 88.33098, 89.6737, 90.91021, 92.39658, 93.70444, 
    94.64077, 90.24769, 91.16688, 92.18113, 93.24791, 94.44572, 96.01465, 
    96.83998, 97.64594, 97.61369, 98.66756, 99.37035, 99.61396,
  83.55575, 85.92578, 88.21295, 90.00874, 91.13099, 91.95337, 92.70006, 
    93.95708, 92.80424, 95.31013, 97.15382, 97.84219, 97.76138, 98.16874, 
    98.75439, 99.31264, 99.71169, 99.86115, 99.9388, 99.92352,
  81.25372, 83.86654, 85.50689, 87.88873, 90.28744, 92.57439, 93.99472, 
    94.992, 95.35307, 95.8008, 96.0643, 96.38999, 96.86933, 97.88213, 
    98.57286, 98.91142, 99.97285, 99.88389, 99.67047, 99.46679,
  78.83917, 80.91822, 82.83163, 84.94747, 86.78602, 88.56271, 89.74208, 
    90.51863, 87.33533, 87.44574, 87.81642, 88.23525, 89.08076, 90.21331, 
    91.41325, 92.43887, 97.4417, 97.80002, 97.94662, 97.52666,
  94.82971, 89.40077, 89.11103, 88.74803, 87.94189, 88.36953, 88.92978, 
    89.50793, 82.19781, 82.37469, 83.71574, 77.99167, 80.06473, 87.88522, 
    88.76618, 87.77132, 93.94604, 94.74261, 95.19641, 95.12885,
  99.00519, 98.81989, 98.04326, 97.91414, 97.95948, 98.42017, 98.41945, 
    98.20856, 95.34817, 95.09523, 94.30952, 93.95645, 94.10553, 96.66939, 
    97.10181, 88.49584, 96.5448, 95.10272, 92.70851, 93.68446,
  97.71663, 97.44809, 97.34927, 97.20062, 96.87726, 96.74217, 96.51619, 
    96.60764, 95.76149, 96.85017, 96.95539, 97.62077, 98.0011, 97.81171, 
    97.58505, 97.17231, 96.93953, 98.34711, 98.97596, 98.72753,
  95.13623, 95.0208, 94.78872, 94.74229, 95.2371, 96.11801, 96.24549, 
    96.57287, 97.10258, 97.40282, 97.30746, 97.38988, 97.32272, 96.53257, 
    96.68906, 96.99647, 97.44928, 98.37415, 98.6228, 98.77359,
  95.1749, 95.25446, 95.36658, 95.40353, 96.50211, 97.21419, 96.77258, 
    96.67493, 96.85016, 97.07955, 96.90733, 96.91724, 96.84129, 96.32203, 
    95.93678, 95.84694, 95.17021, 95.13237, 94.67268, 94.01573,
  93.76662, 93.65955, 93.55228, 93.97215, 94.8518, 93.40412, 85.94259, 
    79.27486, 76.84528, 76.01816, 74.37674, 73.99192, 74.41193, 75.99026, 
    82.06803, 88.64449, 91.21712, 90.22816, 90.76863, 83.60297,
  82.02478, 79.20705, 76.72332, 74.38023, 72.30573, 69.67217, 64.9911, 
    62.30268, 62.1403, 62.3638, 62.14536, 62.3712, 63.15929, 64.31076, 
    66.05291, 67.40738, 68.47811, 69.36456, 69.6653, 67.5464,
  73.08715, 70.78414, 68.54384, 66.98777, 65.30116, 63.70721, 63.00903, 
    63.35164, 64.342, 65.36198, 65.84354, 66.72434, 68.12008, 69.29806, 
    69.87696, 70.6403, 70.34731, 70.24031, 71.21117, 72.79617,
  74.693, 72.27787, 68.94562, 65.9823, 62.90616, 60.96674, 60.90354, 
    62.23541, 63.72224, 65.41039, 67.37131, 69.97499, 72.27907, 73.18038, 
    73.2804, 73.76765, 74.19243, 74.34958, 75.6013, 78.45605,
  72.06964, 70.10696, 64.65933, 59.46721, 57.39639, 58.31934, 60.35738, 
    62.82411, 65.78002, 69.60045, 73.81758, 77.36792, 79.62564, 80.95548, 
    81.50902, 81.48632, 80.63863, 79.29154, 79.82455, 81.63669,
  65.28571, 61.42331, 57.38585, 56.88116, 58.96647, 61.80746, 64.80879, 
    68.42267, 72.15866, 75.72694, 78.95313, 81.9564, 84.12897, 85.59048, 
    85.77937, 84.9611, 82.96798, 80.43719, 78.42764, 77.39595,
  59.93434, 61.3313, 65.14613, 68.3015, 70.92223, 73.30031, 73.38651, 
    70.00507, 67.02206, 66.93287, 69.14425, 73.27285, 77.2766, 80.17863, 
    81.47198, 80.86627, 76.65778, 71.80341, 68.83817, 67.88712,
  67.86378, 73.17168, 76.0937, 76.64691, 76.00099, 72.42905, 65.98078, 
    61.63911, 60.17262, 57.32156, 56.03157, 57.72192, 61.37168, 64.41604, 
    66.4542, 66.77098, 65.27567, 63.82668, 63.56083, 64.4386,
  72.58753, 74.60992, 74.63022, 73.84326, 71.39359, 68.57664, 67.0601, 
    68.20779, 68.48286, 65.45495, 59.89899, 59.97488, 65.75881, 69.31692, 
    69.2757, 69.00771, 69.26047, 69.61372, 70.62437, 72.28876,
  89.96809, 90.15906, 90.71493, 91.28718, 91.62785, 91.91776, 92.71745, 
    93.16669, 91.73727, 92.37442, 92.97276, 93.26537, 93.64071, 93.85204, 
    94.11904, 94.64252, 93.91256, 93.99893, 94.09534, 94.31999,
  85.1158, 86.39758, 87.76208, 89.09888, 90.31291, 91.33238, 92.46342, 
    93.36588, 89.95784, 91.05308, 91.82756, 92.81087, 93.43236, 94.16946, 
    95.34733, 96.08773, 95.08068, 95.89467, 96.89459, 97.72411,
  83.2243, 84.96913, 86.76476, 88.46778, 90.09906, 91.57533, 93.01273, 
    94.09743, 89.3516, 90.21056, 91.62673, 93.13778, 94.17986, 95.58104, 
    96.74451, 97.77769, 97.65915, 98.38472, 98.51648, 98.58967,
  83.99807, 86.01898, 87.6319, 89.24503, 90.80787, 92.17705, 93.24249, 
    93.61642, 91.63387, 93.60515, 95.3684, 96.58596, 97.08095, 97.71061, 
    97.9656, 97.91329, 97.99428, 98.24638, 98.5218, 97.91193,
  81.73453, 82.94801, 84.75771, 86.45647, 88.18287, 89.3878, 90.35136, 
    91.1715, 91.13229, 92.31654, 93.07245, 93.61241, 93.96267, 94.25093, 
    94.3707, 94.48924, 97.65284, 98.12527, 98.46089, 97.59681,
  81.52502, 83.26943, 84.77527, 86.17305, 87.36911, 88.31606, 88.62349, 
    88.59416, 84.84293, 85.29897, 85.76457, 87.09864, 88.50611, 89.75713, 
    90.95892, 92.49658, 98.2957, 99.08614, 99.35757, 98.75723,
  94.12789, 92.07644, 92.33562, 91.99741, 91.23368, 91.12879, 91.31729, 
    91.26303, 83.71767, 85.40928, 87.11419, 80.23, 82.44828, 88.80663, 
    89.9022, 88.11801, 93.303, 94.97079, 96.13844, 96.73497,
  97.78103, 97.83627, 97.65623, 97.06664, 97.22775, 97.72375, 98.37662, 
    98.61763, 95.03325, 94.89096, 93.99583, 94.18608, 95.22114, 98.15991, 
    99.32306, 87.74963, 97.17864, 96.18859, 92.43436, 91.86948,
  98.66531, 98.45119, 98.19391, 98.12972, 98.01772, 97.66002, 97.52949, 
    97.56456, 96.60111, 96.83271, 96.7138, 97.07373, 97.2085, 97.16907, 
    97.67874, 98.22832, 98.42576, 98.80322, 99.005, 98.51038,
  97.82105, 97.28019, 97.30792, 97.42377, 97.43817, 97.42484, 96.82922, 
    96.45273, 96.60254, 96.89478, 97.39455, 97.59484, 97.48067, 96.91296, 
    96.56726, 96.59404, 96.85378, 98.10815, 98.68325, 98.31426,
  96.22511, 96.57211, 96.24015, 96.81547, 97.08661, 97.12953, 97.04643, 
    96.84892, 96.57542, 96.80122, 96.79224, 96.50187, 95.93002, 95.63046, 
    95.46632, 95.55308, 95.35199, 96.31097, 96.84396, 97.57712,
  95.02032, 95.20204, 95.21923, 95.17963, 95.27669, 94.94035, 93.28577, 
    91.6768, 90.15681, 89.46073, 88.50823, 88.44112, 88.19015, 88.78967, 
    92.40214, 93.09899, 92.89092, 93.58162, 94.54745, 93.79881,
  90.30859, 89.94632, 89.13767, 88.02589, 86.32642, 83.25551, 78.7723, 
    74.80079, 72.33775, 70.81233, 69.44589, 69.1961, 70.08909, 71.43599, 
    73.04536, 74.71399, 75.82209, 77.79544, 79.18385, 77.39602,
  81.32109, 79.98638, 77.94798, 75.77444, 73.20747, 70.2383, 68.73551, 
    68.69048, 69.27406, 70.65088, 71.50648, 72.76546, 74.46285, 75.99119, 
    76.62885, 76.59036, 75.40577, 74.57476, 74.26491, 74.35489,
  81.62978, 79.93744, 76.84544, 73.70734, 70.13068, 67.28083, 66.90304, 
    68.28011, 69.75383, 71.58943, 73.61552, 75.86401, 78.03728, 79.47179, 
    80.04943, 80.19865, 79.37127, 78.75881, 78.5974, 79.93369,
  79.83855, 78.18155, 73.2487, 67.80845, 64.71246, 64.73078, 67.02431, 
    69.54002, 71.50209, 74.29035, 77.50314, 79.91391, 81.29193, 81.90332, 
    81.91039, 82.05711, 81.03544, 79.66866, 79.13119, 79.48777,
  73.49921, 68.9416, 63.24607, 61.45179, 62.79889, 65.61633, 68.78905, 
    71.55352, 73.4911, 75.85754, 78.45063, 80.28606, 81.24667, 81.43965, 
    80.5854, 79.4632, 76.75516, 74.10014, 71.87545, 70.05103,
  62.92313, 62.85043, 66.42989, 68.64325, 69.91671, 71.19902, 71.29004, 
    69.08436, 66.83067, 66.75261, 67.8937, 69.65649, 71.42062, 71.75405, 
    71.84883, 71.29756, 67.22771, 62.82701, 60.69414, 60.62553,
  65.47179, 70.83823, 73.38235, 73.00147, 72.30704, 69.5822, 64.19595, 
    61.03735, 60.65143, 58.6284, 57.03741, 57.12055, 57.81227, 58.03138, 
    58.92272, 59.10267, 57.82904, 57.43785, 58.43463, 59.96078,
  65.40292, 66.53486, 67.4348, 67.57095, 66.72198, 64.98051, 62.87617, 
    63.14077, 65.27549, 63.30062, 58.06114, 56.46675, 60.26666, 61.78044, 
    61.75011, 61.63174, 61.6615, 62.31964, 63.69613, 65.23513,
  91.22835, 91.52891, 91.90426, 92.32645, 92.72013, 93.0495, 93.48946, 
    93.85519, 92.3613, 92.75789, 93.07044, 93.37935, 93.67238, 93.99982, 
    94.33788, 94.62806, 93.83258, 93.81764, 94.25726, 94.6286,
  84.32198, 85.3045, 86.32961, 87.30491, 88.37691, 89.44039, 90.4576, 
    91.61155, 88.44921, 89.58254, 90.59374, 91.62606, 92.64285, 93.54321, 
    94.66562, 95.5806, 94.14861, 95.05351, 96.17571, 96.79216,
  84.14957, 85.69971, 87.02478, 88.41084, 89.7412, 91.09847, 92.11122, 
    93.08495, 88.9121, 89.72446, 90.54192, 91.40338, 92.46888, 93.57342, 
    94.55862, 95.33235, 93.93278, 94.55692, 95.02907, 95.68382,
  85.69888, 87.46676, 89.18768, 90.6719, 92.31604, 93.64696, 94.79214, 
    96.01681, 93.76501, 94.40177, 95.15594, 95.82668, 96.46256, 96.78388, 
    96.90022, 97.27876, 97.68348, 97.64367, 97.52276, 97.20686,
  83.26019, 85.33219, 87.44392, 89.16824, 90.79617, 92.13233, 93.12491, 
    94.1566, 93.57332, 93.93491, 94.57185, 95.37153, 96.02441, 96.4966, 
    96.70053, 96.85809, 99.11005, 98.38558, 97.5045, 96.97178,
  83.51756, 84.51206, 84.578, 85.56797, 86.73222, 87.9755, 88.70804, 
    89.17399, 84.90678, 84.68009, 84.614, 84.79279, 85.2931, 85.51572, 
    85.73878, 86.96079, 93.82928, 94.38929, 94.42696, 93.56378,
  92.70278, 90.53497, 90.37027, 90.38954, 90.0672, 90.23486, 90.19421, 
    90.16104, 81.44037, 81.04606, 81.39719, 76.64175, 77.23565, 81.64278, 
    82.62213, 80.76571, 87.18693, 89.16403, 90.54073, 91.45415,
  96.02435, 95.18755, 94.00865, 93.54825, 94.01272, 94.18687, 94.15141, 
    94.06964, 88.97534, 89.05211, 88.39385, 86.61993, 87.89155, 92.45065, 
    94.93445, 82.322, 93.00089, 92.34523, 89.18336, 90.52516,
  96.27517, 95.91504, 95.32773, 94.80378, 94.27042, 93.82578, 93.08898, 
    92.467, 90.85963, 91.07164, 91.0445, 91.09605, 91.98411, 92.50045, 
    93.64713, 94.58318, 95.10674, 96.27628, 95.13901, 95.40903,
  95.10927, 95.06757, 95.4446, 95.56143, 95.76157, 95.20446, 94.60815, 
    93.91383, 93.70384, 93.45914, 93.76832, 93.6042, 93.49659, 93.60081, 
    94.02419, 94.11789, 94.08751, 94.48578, 95.14511, 95.09082,
  94.43353, 94.24761, 94.6473, 94.95407, 95.26637, 94.87921, 94.25951, 
    93.91366, 94.18681, 93.71813, 93.21169, 93.01386, 93.02168, 93.49355, 
    93.89482, 93.89176, 93.0598, 92.8578, 93.30416, 93.8365,
  94.23291, 93.7069, 93.16791, 92.63239, 92.48586, 92.89615, 92.47404, 
    91.19368, 90.08318, 88.06808, 86.04807, 84.7235, 83.80251, 84.28851, 
    85.4758, 87.02997, 87.44542, 88.07337, 89.05791, 90.11639,
  91.77057, 90.32721, 88.80693, 87.55973, 86.35587, 83.7037, 79.508, 
    76.56675, 74.28225, 71.57569, 68.6723, 66.29622, 65.39713, 66.09927, 
    68.3849, 70.94612, 73.17194, 75.39292, 77.0697, 76.99127,
  87.19802, 85.54823, 83.43486, 80.80279, 77.78146, 74.88395, 73.17439, 
    72.45867, 72.11951, 71.76836, 71.10268, 70.86102, 71.69516, 73.33527, 
    74.74741, 75.44687, 74.82057, 74.71159, 75.57297, 76.62046,
  86.9715, 84.56121, 80.65832, 77.14108, 73.07304, 70.11197, 69.23022, 
    70.02097, 71.31416, 72.79099, 74.59866, 76.72959, 78.7088, 79.61921, 
    79.66076, 79.50486, 78.5895, 78.00864, 78.58263, 80.80433,
  83.43156, 81.43723, 76.61904, 71.59091, 68.30677, 67.76372, 69.08311, 
    71.3666, 73.68257, 76.21642, 79.16014, 81.86538, 83.54108, 83.76995, 
    83.37154, 83.22461, 82.29125, 80.60918, 80.24697, 81.37912,
  79.11787, 75.11327, 69.73141, 67.21833, 67.92039, 69.60406, 71.65412, 
    73.81704, 75.80035, 77.98751, 79.85872, 81.76134, 83.15455, 83.77686, 
    84.0577, 83.663, 81.54706, 78.90471, 76.88433, 75.31091,
  70.98434, 69.48456, 71.73927, 73.11094, 74.49874, 75.82857, 75.27575, 
    71.9697, 68.6705, 67.17562, 67.62216, 69.78057, 73.28654, 76.28865, 
    78.11987, 78.12723, 74.67474, 69.7943, 66.2882, 64.48853,
  71.02026, 74.12534, 76.0715, 75.74083, 74.51241, 71.77665, 66.88206, 
    62.82467, 59.63378, 55.43921, 54.12319, 55.94824, 59.3431, 61.47651, 
    62.61919, 62.52587, 60.90301, 59.7467, 59.68172, 60.82912,
  69.75559, 69.48951, 69.63219, 69.80999, 68.3994, 66.41119, 63.33255, 
    60.30617, 60.73796, 57.96996, 55.42238, 56.17302, 61.05106, 62.70873, 
    61.66591, 61.29263, 61.6291, 62.44217, 63.74585, 66.12946,
  91.91817, 92.1753, 92.3112, 92.4333, 92.58778, 92.81447, 93.08449, 
    93.35062, 91.80905, 91.99504, 92.22836, 92.48469, 92.58153, 92.70367, 
    92.91091, 93.14479, 92.31715, 92.54077, 92.66181, 92.73782,
  86.24166, 86.97887, 87.7792, 88.51237, 89.30659, 90.18863, 90.96458, 
    91.83149, 88.34736, 89.0624, 89.80249, 90.56976, 91.38797, 92.14223, 
    92.83375, 93.59395, 91.58875, 92.237, 92.69824, 93.23388,
  83.45387, 84.60576, 85.99773, 87.53622, 89.00977, 90.52225, 91.81526, 
    93.11623, 88.77076, 89.80863, 90.82191, 91.90571, 92.72597, 93.65811, 
    94.43398, 95.12107, 93.26325, 93.89391, 94.46807, 94.99685,
  83.58656, 85.06249, 86.35942, 88.02857, 89.7339, 91.36799, 92.96249, 
    94.8189, 92.25152, 93.27708, 94.11802, 94.33737, 94.65162, 95.01426, 
    95.23357, 95.43066, 96.19344, 95.94753, 95.8487, 95.40548,
  82.24181, 84.14627, 85.97177, 87.8778, 89.43796, 91.14991, 92.49356, 
    93.71217, 92.68405, 93.26865, 93.44203, 93.71092, 93.83102, 94.0048, 
    94.06339, 93.79872, 97.76655, 97.65988, 97.24366, 96.40057,
  82.74071, 85.02032, 86.87373, 88.09276, 89.17245, 89.8027, 90.13021, 
    90.33139, 85.91198, 86.03214, 86.39819, 87.04992, 87.76042, 88.74734, 
    89.79562, 91.1243, 97.26793, 97.69109, 97.86907, 97.45387,
  88.54578, 87.30544, 87.25079, 87.89252, 88.18465, 88.17533, 87.79857, 
    87.34749, 79.33959, 79.91103, 79.66999, 78.04173, 79.05, 83.61814, 
    84.39821, 85.04257, 92.34368, 94.31476, 95.60213, 96.27172,
  91.10552, 91.5318, 91.91953, 91.88432, 91.61529, 91.33934, 91.05523, 
    90.89688, 85.96338, 86.07797, 83.05507, 83.99339, 85.35159, 90.25478, 
    90.03545, 77.37002, 88.04517, 93.29739, 92.89428, 94.43005,
  94.94595, 95.22337, 95.2401, 95.01038, 94.66116, 94.21768, 93.70343, 
    93.09791, 91.0455, 91.17506, 91.48244, 90.83386, 90.03716, 89.53082, 
    89.89446, 90.91457, 90.86484, 91.84815, 91.14241, 93.21554,
  97.14388, 97.46133, 97.52761, 97.47862, 97.73273, 97.36008, 96.91904, 
    96.76087, 96.77469, 96.59953, 96.67117, 96.71708, 96.38613, 95.326, 
    93.93125, 93.89989, 93.88195, 94.02693, 94.29345, 94.36948,
  96.79172, 97.27707, 97.30074, 97.05861, 97.06621, 97.02863, 96.93056, 
    97.03901, 97.34903, 97.09512, 97.03434, 97.29715, 97.50568, 97.47587, 
    96.45058, 96.06673, 96.05328, 95.9228, 95.77122, 95.72007,
  95.05836, 95.20229, 94.7211, 94.41302, 93.98306, 93.19019, 92.51344, 
    91.98919, 91.29247, 90.73058, 89.96471, 90.12168, 91.71012, 93.25563, 
    93.224, 91.36003, 91.20042, 91.82768, 90.95815, 90.51277,
  91.7224, 89.59755, 87.47646, 86.02547, 85.11874, 83.36525, 80.5946, 
    79.95129, 80.2313, 79.82845, 79.33048, 80.21992, 82.10534, 83.86208, 
    84.22647, 83.14131, 81.92301, 81.70592, 81.92039, 81.26216,
  91.90488, 89.76814, 86.07068, 82.68719, 79.74541, 77.19193, 75.96572, 
    76.08807, 76.91937, 78.04131, 78.4928, 79.68465, 81.6516, 83.32336, 
    84.17161, 83.2626, 81.18312, 79.81155, 80.34005, 81.39557,
  88.87624, 86.87465, 82.3545, 77.60839, 73.37327, 71.01565, 71.206, 
    73.06464, 75.89104, 77.78822, 79.35813, 81.36508, 83.68845, 85.34801, 
    85.51057, 84.62672, 82.5945, 81.20314, 80.69298, 81.90855,
  82.56483, 80.9309, 75.2171, 69.04568, 65.96907, 66.55416, 70.04605, 
    74.10661, 77.7887, 80.52696, 82.62484, 84.95423, 87.11452, 88.18942, 
    87.60461, 86.58139, 84.73788, 82.79983, 81.53172, 81.3145,
  74.14912, 70.36305, 65.20955, 63.52248, 65.13507, 68.48318, 72.4311, 
    75.64905, 77.9873, 79.55049, 80.8737, 82.62867, 84.44594, 85.40325, 
    85.71329, 85.41826, 83.13454, 80.86852, 78.99407, 77.31986,
  67.19765, 66.3288, 68.5973, 70.51056, 72.91965, 74.8997, 74.92889, 
    71.96973, 68.20506, 67.1697, 68.09977, 70.88065, 74.46168, 77.27324, 
    80.0017, 80.37282, 77.8334, 74.33208, 72.05119, 70.89472,
  71.83863, 75.07059, 77.05853, 76.29211, 75.18029, 72.63929, 68.80449, 
    65.41692, 61.46516, 58.69772, 57.91452, 59.68964, 64.14354, 68.38145, 
    70.26147, 70.6349, 69.65572, 68.58455, 67.97749, 68.5546,
  75.23919, 74.31561, 72.70142, 70.7337, 69.03269, 67.07004, 65.33653, 
    63.66944, 64.60283, 64.98732, 63.94138, 64.11446, 69.08071, 72.6065, 
    71.9184, 70.68056, 69.97124, 70.12459, 70.91595, 71.97805,
  93.03572, 93.17818, 93.07803, 93.20129, 93.35974, 93.38083, 93.53302, 
    93.72282, 92.26048, 92.57698, 92.84275, 93.41949, 93.84661, 94.1688, 
    94.27666, 94.33641, 93.36643, 93.59779, 93.58037, 93.58857,
  87.17156, 87.98553, 88.50614, 89.00391, 89.47346, 90.09238, 90.69989, 
    91.16663, 87.72911, 88.34229, 89.01591, 89.60275, 89.98563, 90.52453, 
    91.04148, 91.3884, 89.0812, 89.56472, 89.95954, 90.38289,
  83.74214, 84.85846, 86.01733, 87.1892, 88.29929, 89.22572, 89.70461, 
    90.64513, 86.13013, 86.91822, 87.43073, 88.52036, 89.30064, 90.13819, 
    90.85973, 91.61768, 89.53977, 89.91845, 90.42123, 90.89275,
  82.30401, 83.83867, 84.70319, 85.07378, 85.68385, 86.08645, 86.57487, 
    87.15329, 84.11214, 84.96664, 85.84905, 86.6157, 87.68911, 88.60311, 
    89.35109, 90.16465, 91.04706, 90.92582, 90.92285, 90.65399,
  80.32497, 82.47836, 84.33932, 85.66091, 86.80232, 87.77689, 88.59954, 
    89.67031, 88.39588, 88.82681, 89.19852, 89.30243, 89.44788, 89.55249, 
    89.28646, 88.71935, 93.25339, 92.80374, 92.3947, 91.66429,
  80.81848, 83.23454, 85.29358, 87.15211, 87.80119, 88.77476, 89.70412, 
    89.89877, 85.59506, 86.03867, 86.63637, 87.33739, 88.06367, 89.1898, 
    90.17881, 90.72044, 96.5012, 96.46308, 96.4081, 95.84963,
  86.83652, 84.41356, 83.70734, 84.28732, 84.53998, 84.757, 84.65198, 
    84.68118, 77.06798, 76.59726, 75.03759, 77.74955, 79.76186, 84.65909, 
    86.23949, 88.45, 95.14108, 96.77238, 97.37347, 97.65273,
  89.71319, 89.80878, 89.97436, 90.27372, 90.45741, 90.32302, 90.48255, 
    90.39806, 83.45234, 80.56636, 76.36421, 82.43346, 84.51976, 90.35268, 
    84.47293, 79.21237, 79.97634, 94.15541, 92.95548, 94.49334,
  92.75242, 92.59995, 92.54846, 93.17971, 93.61966, 93.67027, 93.57723, 
    93.24665, 89.91059, 88.75574, 88.26729, 87.83854, 87.6041, 88.04456, 
    89.43537, 90.50182, 91.4254, 90.62619, 92.68021, 95.37431,
  92.73845, 93.37518, 94.55936, 95.56993, 95.52206, 94.60944, 94.16314, 
    93.83635, 94.19069, 93.17024, 91.80686, 90.8866, 90.52559, 90.22661, 
    90.22415, 90.65829, 91.68185, 92.86227, 93.33411, 93.66043,
  88.46736, 89.46173, 90.80144, 91.85989, 91.92009, 91.49998, 91.66103, 
    92.07775, 92.90208, 92.11379, 90.97099, 89.80291, 89.49657, 89.4448, 
    89.2961, 89.00839, 88.92309, 89.15536, 89.57014, 90.1797,
  84.81236, 85.77599, 86.75153, 87.88931, 88.69614, 89.03106, 89.11893, 
    89.83617, 90.65471, 90.58871, 89.6525, 88.8248, 88.52641, 88.3697, 
    88.20097, 87.93677, 88.03803, 88.26362, 88.28915, 88.11842,
  88.97031, 89.06528, 88.6657, 88.09039, 87.25834, 85.7926, 83.78144, 
    83.45614, 85.06004, 85.85907, 85.02396, 84.02224, 84.49271, 85.96043, 
    87.28581, 87.59615, 87.41074, 87.10183, 87.20812, 87.32923,
  89.69324, 88.3159, 85.71443, 82.68856, 79.85279, 77.61374, 76.71938, 
    77.14848, 78.28808, 79.94706, 81.1678, 82.27078, 84.08876, 85.99454, 
    87.75903, 88.64365, 87.81761, 87.32012, 87.31942, 87.90106,
  88.8084, 86.90608, 82.86219, 78.6748, 74.24994, 71.32151, 70.83752, 
    72.34718, 74.79339, 77.83905, 80.68529, 83.27451, 85.63631, 87.38405, 
    88.29357, 88.52907, 88.28749, 87.81944, 88.27152, 89.80609,
  84.78685, 82.97536, 77.87247, 72.80954, 70.05477, 69.70261, 71.55586, 
    74.66766, 78.0808, 81.43752, 83.89613, 85.6332, 86.88802, 88.07706, 
    88.48154, 88.58199, 88.57477, 87.96056, 87.58159, 87.90468,
  78.77505, 75.20041, 70.71725, 69.59953, 71.42615, 73.61833, 75.87695, 
    78.29902, 80.22515, 81.52885, 82.69379, 83.85344, 84.59699, 85.40249, 
    85.07623, 84.85587, 83.88961, 82.48152, 81.06894, 79.88236,
  74.05064, 73.79861, 76.08863, 77.99157, 79.31879, 79.66553, 78.17411, 
    75.24071, 71.1261, 69.53804, 70.80364, 73.50418, 75.93468, 77.05521, 
    77.27051, 77.12061, 74.8025, 71.97951, 70.80782, 71.18426,
  79.24635, 82.76532, 83.30587, 81.44402, 79.52573, 76.76073, 72.61305, 
    67.26413, 61.14869, 58.55228, 58.91964, 61.19049, 64.2411, 67.15579, 
    69.1943, 69.81534, 68.98713, 68.41048, 69.25359, 71.32464,
  78.32772, 77.9363, 75.10796, 73.49274, 72.40834, 70.31206, 66.65681, 
    59.49401, 58.68624, 59.91509, 60.50298, 61.85524, 68.00053, 72.92605, 
    74.21884, 74.40737, 73.72869, 73.77547, 74.79834, 76.22893,
  92.09266, 92.37874, 92.61239, 92.87888, 93.16799, 93.46854, 93.75138, 
    94.03291, 92.54502, 92.71645, 93.015, 93.26021, 93.49384, 93.91045, 
    94.25148, 94.38291, 93.7177, 93.78616, 93.74122, 93.62508,
  87.02024, 87.50018, 88.27194, 89.04002, 89.69774, 90.86107, 91.85827, 
    92.62337, 89.35551, 90.03667, 90.56727, 91.11555, 91.69335, 92.33654, 
    93.10432, 93.75599, 92.0074, 92.44286, 92.78152, 93.12635,
  82.97328, 84.09554, 84.82106, 85.74249, 86.61486, 87.46594, 89.14606, 
    90.69543, 87.25216, 88.72365, 89.95661, 90.59101, 91.11993, 91.71912, 
    92.56758, 93.17237, 91.35978, 91.57586, 91.38652, 91.42831,
  83.87892, 85.05746, 86.02435, 86.66299, 87.42369, 88.01917, 88.98538, 
    89.6878, 86.81928, 87.21138, 87.62003, 87.73106, 88.55795, 88.92237, 
    89.34732, 89.65034, 90.47437, 90.43933, 90.70178, 90.79314,
  83.85297, 85.98877, 87.57653, 88.92605, 89.62437, 90.02942, 90.26662, 
    90.87954, 89.42888, 89.82721, 89.94859, 89.39673, 89.33012, 88.8396, 
    88.80294, 88.59731, 93.01898, 92.82733, 92.42233, 91.97584,
  83.39753, 85.70737, 87.71297, 88.75329, 89.55901, 89.55054, 89.70348, 
    90.03745, 86.05724, 86.4035, 86.95789, 87.35156, 87.83746, 88.65073, 
    89.83241, 90.85579, 97.17086, 97.27329, 97.29985, 96.82184,
  88.3615, 85.73872, 84.95748, 85.04754, 84.9671, 84.83407, 84.35245, 
    83.62174, 75.51868, 74.45661, 73.69099, 74.93123, 76.40596, 80.4413, 
    80.06749, 83.82816, 92.02511, 94.47326, 95.70553, 95.92178,
  93.06187, 93.19019, 92.74737, 92.0376, 91.41456, 90.65072, 89.20811, 
    86.79054, 77.53137, 74.75082, 73.3282, 76.91505, 75.81914, 77.04137, 
    67.01234, 70.37905, 73.3315, 90.69579, 91.3021, 92.85958,
  84.87269, 85.38031, 85.33826, 85.31688, 85.8419, 87.19706, 88.90544, 
    89.80481, 86.76443, 85.22227, 83.88287, 82.63313, 82.47033, 82.9679, 
    84.298, 85.71014, 87.89816, 87.63682, 90.95826, 93.89898,
  82.09962, 82.80048, 82.91769, 82.69578, 81.81839, 81.49507, 81.99633, 
    83.30586, 84.40349, 83.97013, 83.22975, 83.61124, 85.15224, 86.689, 
    87.79648, 88.54947, 89.96033, 92.15585, 94.05758, 95.02911,
  83.10207, 84.04843, 84.64211, 84.42923, 83.61931, 82.54053, 81.73926, 
    81.84462, 82.68686, 83.14606, 82.97873, 83.21439, 84.41735, 85.93771, 
    87.33829, 88.31007, 89.42461, 90.5059, 91.72177, 93.28294,
  86.18393, 86.72665, 87.55399, 88.32511, 88.1889, 87.44352, 86.01331, 
    85.06368, 84.77199, 84.68651, 84.89946, 85.31667, 86.2345, 87.19603, 
    88.08532, 88.87093, 90.31078, 91.46145, 92.25913, 93.19031,
  88.86063, 88.56728, 88.68649, 89.155, 88.52061, 86.39948, 84.01324, 
    83.16959, 84.17957, 85.19028, 85.30947, 85.10999, 85.73589, 87.28619, 
    88.42604, 89.06159, 89.9308, 91.05173, 92.1346, 92.82572,
  89.81201, 88.19961, 86.03564, 83.25319, 80.29327, 78.33257, 77.86559, 
    78.75013, 80.54739, 82.23273, 83.25383, 84.41883, 85.74661, 87.51855, 
    89.28563, 89.86731, 89.60383, 89.59972, 90.73492, 92.19923,
  88.48553, 86.08518, 82.45104, 78.76474, 74.741, 72.28807, 72.44984, 
    74.17461, 77.10062, 80.31071, 83.35577, 86.25999, 88.61727, 90.33535, 
    90.74104, 89.93532, 89.02248, 88.89837, 90.29106, 92.50269,
  85.81116, 84.0096, 79.21758, 74.03741, 70.93717, 70.92621, 72.95031, 
    75.99955, 79.87437, 83.84888, 87.25101, 89.54452, 91.02991, 91.66874, 
    91.19263, 90.43174, 89.47283, 89.08804, 89.40852, 90.72321,
  81.64825, 78.51588, 73.63541, 71.14014, 72.38353, 74.5798, 76.82985, 
    79.40304, 82.14717, 84.66114, 86.52576, 87.82308, 88.44505, 88.66312, 
    88.67861, 88.51154, 87.67212, 86.45979, 85.73508, 85.81011,
  76.40799, 74.64326, 74.80235, 75.96683, 77.8071, 79.01524, 78.74644, 
    76.45221, 73.17555, 72.47295, 74.50392, 78.12489, 81.09581, 82.94003, 
    84.92853, 85.36095, 83.29577, 80.43576, 78.99051, 78.84122,
  76.13998, 77.53171, 77.81718, 76.70561, 76.0808, 73.94486, 69.98415, 
    65.09245, 60.4961, 59.36329, 61.0253, 64.53312, 69.50502, 74.37361, 
    77.58986, 78.24058, 76.8185, 75.07291, 74.80775, 76.19957,
  72.69376, 71.56331, 69.71387, 67.95688, 66.70872, 64.99695, 62.56661, 
    58.72014, 59.34329, 61.16765, 63.28808, 64.89376, 69.13304, 73.01115, 
    74.84834, 75.72343, 75.3675, 75.39042, 77.1305, 79.41043,
  91.72614, 91.97892, 92.24584, 92.6017, 92.90726, 93.23003, 93.60563, 
    93.99317, 92.49765, 92.76342, 93.0871, 93.42917, 93.6701, 94.0365, 
    94.2623, 94.41351, 93.55587, 93.63628, 93.89251, 94.03265,
  84.14518, 85.07586, 86.1155, 87.14783, 88.25138, 89.43262, 90.60426, 
    91.707, 88.46263, 89.59267, 90.58944, 91.57991, 92.47266, 93.54031, 
    94.40291, 95.18852, 93.3056, 93.994, 94.62192, 95.14048,
  83.44198, 84.93168, 86.54518, 88.23358, 89.89073, 91.60903, 92.98181, 
    94.19492, 89.77947, 90.99497, 91.84503, 92.91472, 93.81614, 94.66514, 
    95.4581, 96.14622, 94.50372, 95.13116, 95.6834, 96.32315,
  85.90291, 87.40739, 89.07933, 90.7915, 92.36508, 93.66728, 94.8648, 
    95.88739, 93.85136, 94.75296, 95.50141, 96.02695, 96.40417, 96.55314, 
    96.57938, 96.67484, 97.44611, 97.25126, 97.20976, 97.3756,
  86.30454, 88.66948, 90.77248, 92.64782, 93.88834, 94.8798, 95.82591, 
    96.47375, 95.53883, 95.95706, 96.28616, 96.28149, 96.19474, 96.35268, 
    96.24451, 96.07043, 98.60696, 98.25945, 97.69043, 97.0032,
  86.34664, 88.49377, 90.76771, 92.03596, 93.0609, 93.61858, 94.13875, 
    94.30449, 90.0348, 90.24645, 90.7345, 91.1532, 91.43727, 92.34852, 
    93.28825, 94.06742, 98.7078, 98.89421, 98.62544, 97.92306,
  91.76129, 90.27886, 89.54936, 90.19298, 90.01091, 89.42776, 88.91763, 
    88.611, 80.4463, 80.19552, 80.11096, 80.78912, 81.60088, 86.43227, 
    89.33938, 87.27235, 93.84152, 95.8061, 96.80018, 96.7455,
  80.19403, 77.10677, 73.64381, 72.0275, 71.45689, 71.68865, 71.7021, 
    71.62277, 65.87908, 64.67995, 63.78658, 66.84795, 66.1896, 70.10239, 
    70.99362, 75.59287, 84.60676, 88.55972, 87.78676, 89.05531,
  71.63784, 70.08855, 69.5598, 70.25185, 71.41782, 73.34878, 74.83501, 
    75.78947, 73.89905, 74.42846, 74.98672, 75.79089, 77.3736, 79.87261, 
    80.96358, 81.11364, 79.36723, 75.8231, 80.34511, 83.75332,
  77.03259, 77.26087, 76.77525, 76.08031, 75.87844, 76.51199, 77.79214, 
    78.95224, 78.76668, 78.19334, 78.91817, 80.24926, 81.57702, 82.95593, 
    84.30759, 85.43809, 86.62601, 86.86282, 86.32402, 85.20561,
  81.90553, 82.51287, 82.47397, 81.2606, 80.12249, 79.72118, 79.71456, 
    80.27686, 80.64936, 80.23322, 80.25098, 80.33074, 81.10367, 82.28625, 
    83.96735, 85.39771, 86.63801, 87.40573, 88.09508, 88.66438,
  86.2456, 86.40807, 86.81409, 86.70692, 86.42616, 86.20202, 85.46281, 
    85.29221, 84.81882, 84.15075, 83.87453, 84.28586, 84.89616, 85.29898, 
    85.48932, 85.89087, 87.43224, 89.85146, 90.72992, 90.54893,
  89.1325, 88.22382, 88.20148, 88.73246, 88.5392, 87.10438, 85.50205, 
    85.31989, 85.6103, 85.44967, 85.30218, 85.7251, 86.42917, 87.38668, 
    87.72176, 87.53499, 87.84741, 89.09399, 90.04604, 90.83098,
  91.29373, 89.9676, 88.47495, 86.55795, 84.10509, 82.69894, 82.88194, 
    83.93911, 85.24743, 86.28143, 86.54827, 86.85078, 87.77343, 89.28324, 
    90.19785, 89.75495, 88.09054, 87.51006, 88.09782, 88.97469,
  89.86649, 88.2246, 85.18929, 83.0657, 81.3436, 80.54247, 81.31598, 
    83.07146, 84.58733, 86.02483, 87.09673, 88.01353, 88.88243, 89.62682, 
    89.95633, 89.18774, 87.35757, 85.95741, 86.41151, 88.04488,
  86.339, 84.88105, 81.51199, 79.68417, 78.88383, 79.35464, 81.17761, 
    83.1702, 84.97621, 87.00625, 88.49455, 89.38412, 90.08819, 90.34418, 
    89.62489, 88.38779, 86.65417, 85.43839, 85.68197, 86.08061,
  80.83109, 79.23737, 77.70421, 77.78459, 78.49709, 79.57594, 80.43286, 
    81.83361, 83.56165, 84.89755, 86.17075, 87.24276, 87.90272, 87.90722, 
    86.92007, 85.80197, 83.73489, 81.9249, 81.24812, 80.89931,
  75.77617, 75.58641, 77.0136, 78.24151, 78.0391, 77.39792, 76.43443, 
    75.66836, 74.04256, 73.23172, 74.68794, 77.94301, 81.02079, 82.66119, 
    82.43949, 81.05273, 78.17992, 75.69452, 75.13483, 74.97328,
  72.17251, 74.30869, 74.50819, 73.38627, 71.6301, 71.07693, 69.62086, 
    66.7551, 64.47157, 63.52911, 63.78706, 65.79415, 69.61604, 72.12495, 
    73.40547, 73.1663, 72.57866, 71.77567, 71.98804, 72.67963,
  66.01498, 65.5641, 63.7215, 63.7728, 65.77634, 67.18826, 67.42655, 
    64.69852, 65.98106, 67.45634, 67.5254, 67.70526, 70.16753, 71.7878, 
    72.78249, 73.43069, 73.33083, 73.33017, 73.91627, 73.78754,
  92.7289, 93.1573, 93.54835, 94.08183, 94.45391, 94.84051, 95.25007, 
    95.63009, 94.73144, 95.07844, 95.47897, 95.81799, 96.03333, 96.26595, 
    96.43076, 96.65799, 96.24045, 96.44221, 96.74995, 96.62806,
  88.14227, 89.29109, 90.46381, 91.55473, 92.56074, 93.45291, 94.2736, 
    95.17516, 92.1431, 92.81657, 93.50533, 94.24451, 95.28857, 96.21684, 
    96.95387, 97.57932, 96.40977, 97.20378, 97.74783, 98.13219,
  88.14897, 89.59606, 90.8746, 92.18648, 93.4766, 94.69495, 95.85283, 
    96.89256, 92.81134, 93.77935, 94.74272, 95.78279, 96.57649, 97.25861, 
    98.08129, 98.70869, 97.46019, 97.77924, 97.98026, 98.51221,
  87.39945, 89.04401, 90.70658, 92.34492, 93.93926, 95.42852, 96.43814, 
    97.15221, 94.52446, 95.37478, 96.17605, 96.82298, 97.44414, 98.06287, 
    98.46099, 98.67272, 99.01943, 97.60178, 97.11073, 97.50469,
  86.46487, 88.17768, 90.33053, 92.37748, 93.87351, 94.97795, 95.97858, 
    96.65021, 95.71638, 95.82104, 95.57257, 94.9843, 94.56375, 94.51633, 
    94.51193, 94.63573, 97.3384, 96.74677, 96.6872, 96.67126,
  86.14116, 88.17406, 90.20102, 92.0609, 93.16382, 93.76161, 94.05056, 
    94.32043, 89.20064, 88.25187, 86.80096, 86.14659, 86.56003, 87.01359, 
    87.32991, 87.48611, 93.7278, 94.35239, 94.62696, 94.00191,
  93.18294, 92.58247, 92.65812, 92.96688, 92.91366, 93.07026, 92.12991, 
    91.01332, 82.99873, 82.56676, 81.44022, 76.54862, 77.71646, 83.14697, 
    86.34957, 81.52479, 88.51782, 91.09167, 93.06666, 93.33993,
  75.1904, 71.68581, 69.46727, 68.24815, 67.95087, 68.70954, 67.49162, 
    65.69518, 59.46147, 58.31851, 59.05737, 65.77574, 71.91098, 83.52595, 
    89.04636, 89.99678, 91.75639, 90.83635, 86.90574, 86.33804,
  70.90353, 70.48632, 70.57195, 70.59414, 70.4999, 70.81147, 71.25254, 
    71.67159, 70.37982, 70.57768, 70.40791, 70.73579, 71.55083, 73.8223, 
    74.18034, 74.69206, 77.7923, 83.56129, 87.65398, 89.59861,
  77.72495, 77.64016, 77.70279, 77.73128, 77.63654, 77.45772, 77.3634, 
    77.43354, 78.18114, 78.77745, 79.69411, 80.72012, 81.15813, 81.53223, 
    81.17523, 80.60073, 79.89496, 79.94285, 79.64116, 79.12093,
  82.40411, 82.0882, 81.72245, 81.62374, 81.83842, 81.88451, 81.8376, 
    82.16739, 83.12712, 83.13606, 83.4146, 84.05341, 84.88135, 85.5474, 
    86.09451, 86.82574, 87.412, 87.84286, 87.98222, 88.07838,
  85.29477, 84.82441, 84.78718, 85.6182, 86.59268, 86.95855, 86.48321, 
    86.51676, 87.31081, 86.92317, 86.42233, 86.44984, 87.18022, 88.24606, 
    89.04674, 89.22823, 88.82217, 89.56557, 90.11314, 89.43811,
  85.51265, 85.32461, 85.9403, 86.54429, 86.44884, 85.08876, 83.43629, 
    82.81059, 83.38242, 83.3542, 83.21011, 83.47954, 84.64256, 86.36319, 
    87.7826, 88.19127, 87.60859, 88.08943, 88.68541, 87.59548,
  86.35654, 85.58758, 84.49693, 82.50793, 80.06528, 78.17739, 77.27887, 
    77.65334, 79.18013, 80.81451, 81.74583, 82.97023, 84.48615, 86.38699, 
    87.84322, 88.03423, 87.01444, 86.49339, 86.68327, 86.5595,
  85.99264, 85.06941, 82.7449, 80.04942, 77.18018, 75.32719, 75.44117, 
    77.20317, 79.92599, 82.01187, 83.78746, 85.64829, 87.18235, 88.00639, 
    88.35136, 87.63506, 86.07841, 84.65396, 85.02084, 86.1767,
  82.8708, 81.88372, 78.25472, 74.86462, 73.17766, 73.60953, 75.5573, 
    78.22768, 81.11987, 83.40513, 85.68612, 87.24898, 87.85596, 87.6541, 
    86.5577, 85.45315, 84.62639, 84.40824, 85.23612, 85.8003,
  76.11572, 74.28699, 72.00488, 71.88872, 73.64548, 75.40047, 77.02804, 
    78.56323, 80.01992, 81.2054, 82.89726, 84.36304, 84.71316, 84.41503, 
    83.78284, 83.92426, 83.95953, 83.99019, 84.07111, 83.89619,
  71.48241, 70.74561, 72.35433, 75.00738, 76.70261, 76.47975, 74.78413, 
    71.83713, 68.65202, 68.75716, 72.23263, 75.94894, 79.18945, 80.94232, 
    82.49986, 84.47905, 84.89851, 82.8448, 80.93427, 79.35069,
  71.10316, 73.89064, 76.53503, 76.40215, 73.39511, 70.12331, 66.3209, 
    62.96446, 62.10137, 63.88395, 66.40358, 70.22091, 74.58755, 77.38135, 
    79.12296, 79.29867, 78.41794, 76.23497, 73.816, 72.41816,
  70.03917, 69.58164, 68.34452, 66.38229, 66.23264, 66.1891, 66.68623, 
    66.60573, 69.91621, 74.07331, 73.81617, 73.97363, 76.49303, 78.04353, 
    77.65372, 76.77383, 75.61914, 73.91495, 71.92735, 71.81947,
  92.99148, 93.38159, 93.82012, 94.33382, 94.79841, 95.13759, 95.73686, 
    96.08545, 94.896, 95.34359, 95.90163, 96.01503, 96.49646, 96.50758, 
    96.93884, 96.94193, 96.48019, 96.68491, 96.74319, 97.36211,
  89.47833, 90.88607, 92.24848, 93.69579, 95.23843, 96.45618, 97.27627, 
    98.04473, 95.3, 96.03017, 96.22168, 96.4677, 96.69855, 96.9447, 97.33379, 
    97.67093, 95.61038, 95.94926, 96.43163, 96.92271,
  90.73714, 93.14381, 95.25055, 96.58489, 97.55779, 98.24677, 98.54967, 
    98.8447, 95.62145, 95.9582, 96.21976, 96.93179, 97.49046, 97.95266, 
    98.11625, 98.32435, 97.33636, 97.841, 98.43262, 99.1521,
  89.63442, 92.39142, 95.03806, 96.8643, 97.5985, 97.9479, 98.22198, 98.5115, 
    96.69513, 97.06969, 97.69389, 98.29397, 98.94601, 99.33304, 99.53901, 
    99.71231, 99.91858, 99.91685, 99.81169, 99.65685,
  86.48783, 90.35569, 92.52915, 93.98511, 94.80739, 95.58295, 95.82641, 
    95.61538, 93.52598, 93.11774, 93.42233, 94.1953, 95.32901, 96.67121, 
    97.81027, 98.58317, 99.97215, 100, 99.99611, 99.94057,
  86.87508, 90.16988, 92.64064, 93.42454, 93.51669, 93.50846, 93.38802, 
    93.10145, 88.8437, 88.89963, 89.25941, 89.99405, 90.52409, 90.32795, 
    89.84596, 90.3817, 95.7711, 96.54607, 97.23893, 97.36222,
  98.29879, 96.88589, 96.3633, 96.28941, 96.01233, 95.85963, 95.24767, 
    94.72495, 86.93438, 86.6211, 86.9519, 81.78722, 82.0987, 84.31771, 
    87.93884, 85.52946, 91.17413, 92.94044, 94.49667, 95.36691,
  93.78554, 90.59438, 86.82793, 85.20072, 85.94543, 88.77772, 90.26144, 
    90.22134, 84.17958, 82.85894, 83.52737, 80.12448, 80.61956, 85.40114, 
    91.25476, 91.80544, 93.42714, 91.50433, 91.23431, 91.77765,
  73.63203, 67.14255, 63.53806, 63.13897, 63.45485, 63.51927, 63.69291, 
    63.4581, 61.75826, 62.40147, 64.3262, 69.44565, 76.23885, 82.1163, 
    83.80643, 84.42504, 86.70598, 90.76015, 93.76917, 94.30648,
  71.03206, 71.78105, 72.99789, 73.70122, 73.34026, 72.33054, 71.15786, 
    70.07006, 69.25307, 68.58427, 68.63718, 69.3344, 69.84557, 70.15797, 
    69.96938, 70.24627, 71.31436, 72.75469, 74.67911, 77.13605,
  78.12453, 77.98836, 77.8632, 77.54881, 77.11539, 76.61423, 76.36926, 
    76.08171, 75.77153, 75.42714, 75.35838, 75.50757, 75.82435, 75.8967, 
    75.71997, 75.79306, 76.28555, 76.70612, 77.51298, 78.49121,
  82.01278, 81.7551, 81.48304, 81.61835, 81.84556, 81.45633, 80.70699, 
    81.01472, 81.00084, 80.60494, 79.87412, 79.77531, 80.46571, 81.4369, 
    81.77026, 81.72459, 81.98112, 82.66138, 83.04337, 81.78686,
  84.21192, 83.91651, 83.80417, 84.11613, 83.95065, 82.75063, 81.22007, 
    81.21228, 81.03355, 80.62953, 79.68715, 79.24458, 79.77376, 81.25245, 
    82.78201, 83.37992, 83.00098, 83.33106, 83.57304, 82.75285,
  85.12054, 84.15527, 83.14683, 81.64615, 79.96709, 78.78537, 78.32475, 
    78.6692, 78.89671, 79.39584, 79.61345, 80.11021, 81.15524, 82.81792, 
    84.43388, 84.71048, 83.7061, 83.24312, 83.41142, 83.39447,
  87.29604, 86.12797, 83.79558, 81.52433, 78.7413, 76.32051, 75.84665, 
    77.28436, 78.83002, 80.29754, 81.6159, 83.10711, 84.5929, 85.6211, 
    86.06468, 85.7447, 84.26506, 83.02289, 83.49651, 84.49574,
  85.7327, 84.64523, 81.29393, 78.43938, 76.32657, 75.64949, 76.79267, 
    78.87111, 80.57969, 82.09154, 83.37271, 84.54805, 85.50865, 85.90814, 
    85.1416, 83.95724, 82.09579, 81.16747, 81.8436, 83.05403,
  80.78965, 78.49258, 76.26681, 76.30175, 77.60586, 78.93127, 79.9437, 
    80.47091, 80.67621, 81.0602, 81.75932, 82.7703, 83.31271, 83.14477, 
    81.84224, 80.26047, 77.99124, 76.6957, 76.2996, 76.73602,
  77.62566, 77.20658, 79.32854, 81.97481, 82.80705, 81.55907, 79.16624, 
    74.48483, 69.56812, 68.30215, 69.89416, 72.73569, 74.64589, 74.54435, 
    73.3232, 72.0088, 69.43981, 67.30808, 66.43539, 66.80431,
  76.4373, 79.4134, 81.51705, 80.72845, 78.64883, 76.93772, 73.77604, 
    68.33348, 64.96485, 62.41588, 60.94473, 60.97815, 61.34219, 61.11619, 
    60.06549, 58.56825, 57.08685, 56.91457, 57.9743, 59.75175,
  72.4187, 72.1474, 71.27704, 72.36794, 74.55864, 75.4277, 73.99171, 
    69.17621, 68.59572, 68.20935, 64.27888, 62.02097, 61.58382, 61.42978, 
    60.41274, 58.74488, 56.64424, 56.17491, 57.81411, 61.17122,
  93.72971, 94.03551, 94.43389, 94.75692, 95.23486, 95.43662, 95.82867, 
    96.24335, 94.89697, 95.18201, 95.56387, 95.81216, 96.11404, 96.44719, 
    96.49788, 96.82176, 95.8974, 96.28552, 96.72123, 96.84827,
  86.61088, 88.01867, 89.42487, 90.89743, 92.22617, 93.45229, 94.57592, 
    95.58984, 91.83442, 92.59222, 93.4392, 94.44369, 94.86494, 95.42963, 
    96.22427, 96.64986, 95.15445, 95.84504, 96.42202, 97.01573,
  88.85981, 90.53657, 91.92621, 93.05698, 93.95808, 94.74271, 95.43624, 
    96.0235, 91.35714, 92.21185, 93.06292, 93.66696, 95.3672, 96.7281, 
    97.32455, 97.71213, 97.01571, 97.59209, 98.02304, 98.33675,
  88.84864, 90.9267, 92.52587, 94.11626, 94.80871, 94.90771, 94.56481, 
    95.05518, 92.73986, 93.33976, 94.31722, 94.90302, 95.96869, 97.09246, 
    97.90607, 98.42188, 99.08035, 99.19006, 98.75628, 97.7698,
  86.80632, 88.5857, 89.93571, 90.63291, 89.48568, 87.88619, 88.28513, 
    88.76382, 88.50789, 88.87151, 89.96033, 91.38094, 92.58386, 93.65589, 
    94.34502, 95.28899, 97.922, 98.89149, 98.91284, 98.27467,
  82.39191, 84.53304, 85.93727, 87.09081, 86.93341, 86.19765, 86.24261, 
    86.58118, 82.3757, 82.14922, 82.38621, 82.94489, 84.40987, 86.68294, 
    89.18845, 91.18963, 97.6476, 98.77509, 99.25974, 99.13137,
  94.49702, 90.6898, 89.86106, 90.46116, 89.80382, 88.86613, 87.43515, 
    86.10226, 77.73002, 78.09724, 79.53412, 73.65804, 74.98666, 80.24499, 
    83.47589, 81.46077, 87.81081, 90.10869, 92.19386, 93.3928,
  89.50273, 87.54592, 86.04684, 85.55839, 86.07019, 86.85114, 87.41547, 
    88.10159, 84.23147, 86.14262, 89.45796, 84.66185, 83.42672, 87.28989, 
    90.76624, 92.63701, 93.22452, 91.66343, 89.1031, 91.10976,
  90.92999, 89.11899, 88.45069, 87.39809, 87.97838, 87.62603, 86.89352, 
    87.10899, 86.01675, 88.3881, 91.63838, 93.45891, 92.08976, 90.96973, 
    90.43681, 91.41393, 93.26367, 95.38046, 95.71567, 95.65543,
  80.15085, 77.99427, 76.7924, 75.89832, 74.16212, 73.36053, 73.47568, 
    73.39588, 72.08852, 71.85829, 74.05017, 76.87769, 79.91053, 79.99729, 
    79.11797, 78.74055, 79.43986, 82.78654, 86.38605, 87.82205,
  76.91962, 77.1038, 77.25069, 77.32476, 76.87509, 75.8241, 74.7005, 
    73.67066, 72.31319, 71.58145, 70.91515, 70.44945, 70.27596, 70.26601, 
    69.76395, 69.4837, 69.57767, 69.82037, 70.35172, 70.29267,
  77.661, 78.18739, 78.58044, 78.91357, 79.1022, 78.10476, 76.41315, 
    76.26118, 76.77834, 76.60896, 75.66179, 75.0564, 75.16804, 75.87793, 
    76.41117, 76.04704, 75.67166, 75.65691, 75.33081, 73.60004,
  78.37594, 78.60741, 78.96687, 79.31673, 78.82134, 76.99261, 75.03725, 
    74.85607, 75.63193, 75.68449, 75.04001, 74.48342, 74.4257, 75.6045, 
    78.09108, 79.62678, 79.54363, 79.09273, 78.29303, 76.1933,
  77.89133, 77.01044, 75.87775, 74.52716, 72.73531, 70.92063, 70.14401, 
    70.6374, 71.30305, 71.90122, 72.30972, 72.78746, 73.64633, 75.6529, 
    79.58994, 81.98377, 81.48635, 80.40215, 79.79695, 79.84991,
  79.04986, 77.96844, 75.58145, 72.76558, 69.30787, 66.75317, 65.99226, 
    66.82247, 68.68903, 70.81125, 72.80035, 75.0694, 77.91127, 80.82827, 
    83.35236, 84.53519, 83.80582, 82.43272, 82.307, 83.36151,
  78.61369, 76.9856, 72.85793, 68.26077, 64.9839, 64.03307, 65.15066, 
    67.98197, 71.69209, 75.22868, 78.22675, 80.82264, 82.95004, 84.7879, 
    85.38228, 85.12318, 84.09585, 83.10471, 83.8761, 84.94166,
  76.22778, 73.07869, 69.35329, 67.88725, 68.99717, 70.82835, 73.11674, 
    75.74903, 78.22446, 80.33199, 82.38418, 83.95488, 84.7705, 85.306, 
    85.11682, 84.40217, 83.11152, 81.87775, 81.24982, 80.99374,
  73.84452, 72.28394, 73.99317, 76.73956, 79.19324, 79.88586, 77.5317, 
    72.29091, 67.98129, 68.12842, 71.13874, 74.55568, 77.78831, 79.48026, 
    80.14385, 80.08586, 77.42348, 74.18307, 73.02173, 73.06721,
  73.63855, 76.6207, 79.05457, 79.02032, 77.79808, 73.94193, 67.00645, 
    61.17018, 60.21066, 58.87897, 58.93137, 59.97506, 61.33646, 62.03708, 
    62.69863, 63.60392, 64.0003, 65.2429, 67.18152, 69.03476,
  70.39806, 71.68782, 71.07378, 69.93989, 69.35001, 67.59538, 65.62215, 
    63.93141, 65.27674, 63.95311, 60.06851, 59.02525, 60.88435, 64.10941, 
    65.81861, 66.63889, 68.33271, 70.43531, 72.28477, 73.37875,
  93.64671, 94.05598, 94.47609, 94.51242, 94.45212, 94.68769, 95.05457, 
    95.25493, 93.67635, 93.72635, 94.31325, 94.46198, 94.7226, 94.78752, 
    95.19112, 95.2608, 94.31791, 94.39255, 94.78739, 94.66754,
  89.65529, 90.74836, 91.91697, 92.89857, 93.53438, 94.55206, 94.93401, 
    95.69736, 91.58758, 92.13486, 92.37679, 93.36708, 93.82729, 94.49367, 
    94.81551, 95.41537, 93.40851, 94.17928, 94.66608, 95.34855,
  86.61282, 88.3792, 90.09097, 91.65804, 92.97572, 94.06114, 95.15382, 
    96.06357, 91.73462, 92.97826, 93.89375, 94.72905, 95.02287, 95.93253, 
    96.66759, 97.69312, 97.68056, 98.53715, 99.19547, 99.70373,
  86.36751, 88.52943, 90.64953, 92.47297, 93.51411, 94.47469, 95.72016, 
    96.40972, 94.69509, 94.59147, 93.43809, 94.66803, 96.5032, 97.64626, 
    98.60197, 99.09479, 99.54364, 99.77277, 99.95231, 99.99925,
  82.87292, 84.81871, 86.33745, 87.62495, 88.56259, 88.01833, 88.79974, 
    89.80191, 89.98247, 91.01443, 91.28108, 92.31226, 93.23839, 94.54628, 
    95.75062, 97.13625, 99.20444, 99.67713, 99.7452, 99.07822,
  82.38123, 82.71155, 82.84904, 83.21956, 83.09562, 82.3077, 82.40763, 
    83.12376, 79.7402, 81.18941, 82.44987, 84.66368, 85.7455, 86.71981, 
    88.09573, 90.00997, 96.57462, 97.27665, 97.34451, 96.77862,
  92.53261, 88.19363, 85.38067, 83.72462, 81.66814, 80.31536, 79.72077, 
    79.95586, 72.89447, 74.32348, 77.4297, 72.43382, 74.4905, 81.82894, 
    84.0457, 81.13492, 87.24388, 89.39352, 91.14304, 91.89108,
  97.08171, 95.16993, 92.76344, 90.67206, 89.96401, 90.64304, 91.83529, 
    94.25391, 91.52099, 92.77678, 94.81535, 91.02692, 89.62936, 93.89788, 
    92.9303, 91.81164, 92.64296, 91.11305, 87.79584, 88.74056,
  98.67889, 98.04272, 96.59895, 95.94193, 96.22273, 96.11771, 96.68858, 
    97.3736, 97.06327, 98.39551, 98.7389, 98.57149, 98.49107, 97.32613, 
    95.14423, 94.63239, 96.09977, 97.47442, 97.80214, 97.05959,
  96.98618, 94.65034, 92.22398, 92.7278, 92.98281, 92.86243, 92.95996, 
    93.85134, 94.93194, 96.53144, 98.17088, 98.77944, 98.55646, 98.5482, 
    97.88772, 97.37463, 97.10835, 97.45614, 98.07851, 98.77384,
  83.01666, 81.56857, 78.75431, 76.536, 75.10692, 73.97153, 73.77499, 
    74.86559, 76.52209, 77.19692, 77.88699, 79.40308, 82.16992, 84.35828, 
    83.48967, 81.21072, 81.05755, 83.22154, 83.14905, 81.51738,
  66.95157, 67.28563, 67.13587, 67.44505, 67.43891, 66.90847, 66.28897, 
    67.12601, 68.73547, 69.20729, 69.11932, 69.21804, 70.10564, 71.07471, 
    71.47787, 71.04275, 70.63866, 71.25925, 70.53139, 68.61951,
  71.35865, 70.21389, 69.60371, 69.58196, 69.21909, 67.93578, 66.72469, 
    67.16914, 68.46863, 69.32945, 70.00468, 70.99332, 72.82994, 75.61628, 
    79.52466, 81.86647, 82.50616, 82.57534, 82.00821, 79.86826,
  73.85767, 72.8142, 71.52262, 69.8084, 67.73034, 65.60339, 64.49372, 
    64.96942, 67.12055, 70.09428, 72.78183, 75.60758, 78.41879, 81.33156, 
    84.60886, 86.60928, 86.36523, 85.93711, 85.16256, 83.85181,
  75.61953, 74.85708, 73.2029, 70.90084, 67.02274, 63.72683, 62.79031, 
    64.78535, 68.99979, 72.97313, 76.2082, 79.33366, 82.09197, 84.17397, 
    85.72778, 86.52843, 86.15574, 85.19884, 84.67241, 84.93076,
  75.13121, 73.84025, 70.06603, 65.19676, 61.22583, 60.04469, 62.33815, 
    67.02165, 72.55351, 76.79778, 79.97818, 82.56522, 85.05787, 87.33788, 
    88.03735, 87.64152, 86.42144, 85.2137, 85.21176, 85.34274,
  68.82114, 65.20398, 60.33849, 57.47905, 57.77803, 60.98416, 65.87654, 
    71.43363, 75.98819, 78.95587, 80.83644, 82.51546, 84.83549, 86.79829, 
    87.26402, 87.12022, 85.97598, 84.34417, 82.93956, 81.10789,
  61.68291, 59.48023, 60.2206, 63.23719, 67.0256, 70.34559, 70.37291, 
    67.21758, 64.75401, 65.19872, 67.91457, 72.31242, 76.97902, 80.82691, 
    82.94274, 83.18847, 80.61556, 76.04985, 71.88647, 68.96687,
  61.12665, 63.32415, 66.28885, 69.18752, 69.56549, 66.41309, 60.21794, 
    55.90883, 56.44659, 56.578, 56.76321, 58.48072, 61.71857, 64.62292, 
    66.14228, 66.09158, 64.54202, 62.12258, 61.18162, 61.79814,
  60.57084, 61.47084, 62.07775, 62.5121, 61.50113, 59.43485, 58.44446, 
    61.42545, 61.71103, 59.59251, 53.63789, 54.33769, 59.35477, 63.1613, 
    63.14772, 62.11299, 61.60023, 61.6436, 62.873, 64.95,
  92.46906, 92.65533, 92.89652, 93.38924, 93.74599, 94.1208, 94.46406, 
    94.77744, 93.24382, 93.61447, 93.89458, 94.16271, 94.49475, 94.75928, 
    94.93324, 94.99646, 94.1124, 94.50582, 94.74752, 94.76996,
  85.44726, 86.7691, 88.10397, 89.52422, 90.80333, 91.88545, 92.77533, 
    93.8353, 90.53826, 91.49055, 93.1425, 94.14516, 95.05296, 95.79193, 
    96.38642, 96.64764, 94.96072, 95.59815, 96.1243, 96.47279,
  84.47685, 85.90644, 87.31581, 88.9323, 90.73951, 92.34937, 93.52151, 
    94.43581, 90.36732, 92.523, 94.51615, 95.7461, 96.61171, 97.43674, 
    97.87655, 98.70796, 98.02767, 98.09313, 97.97078, 98.1229,
  83.77087, 85.96499, 87.99674, 89.94136, 92.14854, 94.02409, 95.05857, 
    95.52141, 94.00761, 95.26956, 96.33098, 97.24252, 97.42923, 98.25863, 
    98.8583, 99.72722, 99.92117, 99.28725, 98.52301, 98.13625,
  77.49356, 78.6956, 79.42404, 80.5606, 82.1739, 82.94969, 84.05997, 
    85.42072, 85.72886, 87.11221, 88.32635, 89.5744, 90.88866, 92.25807, 
    93.60825, 94.97401, 97.7389, 98.20255, 98.54131, 98.62502,
  77.87165, 79.12363, 80.97923, 82.91417, 84.72533, 86.18265, 86.76503, 
    86.81076, 81.63461, 82.1003, 83.20142, 84.72913, 86.55308, 88.43545, 
    89.23932, 90.13791, 96.78021, 97.86923, 98.44961, 97.97797,
  93.23658, 87.46267, 88.26495, 88.73966, 88.42339, 88.26445, 88.47377, 
    88.80663, 81.54901, 81.84605, 82.85259, 76.42375, 78.37042, 86.28273, 
    89.06393, 83.3202, 88.53681, 90.22797, 91.64175, 92.01548,
  97.39009, 97.09064, 97.14641, 97.35262, 97.38901, 97.29236, 97.74508, 
    97.92564, 93.70269, 93.998, 95.0431, 91.77088, 92.40113, 95.25706, 
    96.83901, 89.08591, 95.06578, 94.45523, 90.20075, 90.33872,
  99.4864, 99.3409, 98.84968, 98.78441, 98.58266, 98.28791, 97.85995, 
    97.40744, 95.40929, 96.25834, 96.77511, 96.99531, 97.11633, 96.91389, 
    96.2593, 96.5637, 97.33052, 98.40083, 98.59831, 98.40445,
  97.33491, 96.91238, 96.1853, 95.52367, 95.53385, 95.18797, 94.76951, 
    94.26254, 93.93301, 94.89368, 95.6363, 96.0668, 96.41718, 96.63584, 
    97.27202, 97.87407, 98.26603, 98.48637, 98.5992, 98.87265,
  95.79751, 96.03111, 96.27702, 95.99687, 95.29163, 94.42066, 92.70629, 
    91.76328, 90.82865, 90.46668, 90.84836, 91.19216, 91.47442, 91.79884, 
    92.18448, 92.17316, 92.39298, 92.75448, 93.21896, 92.74178,
  88.34765, 87.64189, 87.04655, 84.50876, 81.10733, 74.3058, 68.82692, 
    67.75849, 69.16976, 70.1438, 71.7377, 73.98956, 76.55395, 79.39594, 
    81.47217, 82.0571, 82.1991, 82.38724, 82.02624, 80.74789,
  72.949, 71.63059, 70.59606, 69.50647, 68.65765, 67.57097, 66.94695, 
    67.71823, 69.508, 71.01711, 72.10677, 73.35306, 74.9211, 77.17082, 
    79.74715, 81.54626, 81.77248, 81.5286, 81.39123, 80.20009,
  73.57469, 72.44406, 71.01122, 69.5947, 67.99151, 66.61679, 66.06182, 
    66.81452, 69.10004, 71.26022, 72.6619, 74.46738, 76.90388, 79.41286, 
    81.62605, 83.2546, 83.27071, 83.13461, 83.13335, 82.76216,
  74.43343, 73.34287, 71.63875, 69.20613, 65.29713, 62.20803, 61.41346, 
    62.94527, 66.32952, 69.24154, 72.13495, 75.59301, 78.7777, 80.88163, 
    82.50214, 84.044, 84.66105, 83.9819, 83.58504, 84.14858,
  72.43533, 70.84338, 66.73032, 61.36561, 57.01369, 55.66636, 57.1587, 
    60.78001, 66.0844, 70.78642, 74.90363, 78.1708, 80.64423, 82.68915, 
    84.4777, 84.73186, 83.61091, 82.43195, 82.89045, 83.90265,
  63.68211, 59.62016, 54.9061, 52.51707, 53.12894, 55.35194, 59.2934, 
    64.10414, 69.98523, 74.39243, 77.86761, 80.73233, 83.15685, 85.25098, 
    85.88614, 84.68256, 82.58968, 80.85189, 79.87296, 79.69402,
  54.7021, 53.76855, 55.7305, 58.29206, 61.5443, 64.83125, 66.24121, 
    64.17365, 62.24245, 62.47628, 66.00048, 71.19569, 76.53123, 79.93232, 
    81.80828, 81.23856, 77.68692, 73.37079, 70.98148, 70.45665,
  60.09565, 63.75784, 66.14206, 67.43174, 67.0727, 63.22318, 57.73834, 
    54.70699, 55.1712, 53.98062, 54.0881, 56.5186, 61.05513, 64.60146, 
    66.44014, 67.22374, 66.92986, 66.34594, 66.4712, 66.99677,
  66.18935, 67.30225, 66.549, 64.08141, 60.11318, 55.88155, 55.11483, 
    60.43969, 61.30338, 59.39874, 54.51205, 56.16283, 62.90117, 69.15146, 
    70.78698, 71.53653, 72.68771, 72.979, 73.115, 72.74686,
  91.89491, 92.12323, 92.44369, 92.70435, 92.98618, 93.13318, 93.51932, 
    93.67699, 92.30843, 92.8224, 93.17683, 93.38063, 93.6017, 93.92322, 
    94.21494, 94.27192, 93.53002, 93.68031, 93.70236, 93.67761,
  87.08045, 87.73311, 88.27898, 88.82833, 89.79833, 90.88193, 92.04939, 
    93.15852, 89.7802, 90.44158, 90.86254, 91.76184, 92.1877, 93.09108, 
    93.61987, 94.4933, 93.00451, 93.87434, 94.78695, 96.56996,
  86.57347, 87.17926, 87.925, 88.70908, 89.62112, 90.52332, 91.46152, 
    91.91439, 86.73261, 87.12942, 88.01848, 89.76748, 91.20564, 92.09039, 
    92.96558, 94.10017, 94.09179, 95.77605, 97.09556, 98.29575,
  85.40817, 86.22214, 87.28826, 88.03706, 88.79945, 90.5043, 91.99727, 
    92.72769, 90.43909, 91.64767, 92.91025, 94.44183, 96.74718, 98.62967, 
    99.03271, 97.82977, 97.04924, 96.86734, 97.24192, 97.77924,
  82.38597, 83.04021, 83.35707, 83.06908, 83.99233, 85.09217, 86.76245, 
    88.05067, 88.41999, 89.80721, 91.39365, 92.89558, 93.95396, 94.76693, 
    95.53843, 96.46169, 99.17386, 99.44891, 99.18778, 98.41818,
  79.90095, 80.19803, 80.53106, 81.74171, 82.67239, 83.95, 85.13409, 86.3401, 
    82.85722, 83.48864, 84.33512, 85.24976, 86.1935, 87.37616, 88.66477, 
    90.10486, 96.30755, 97.25281, 97.24182, 97.40324,
  94.02654, 90.63446, 89.37109, 87.34268, 86.04471, 85.48306, 85.40534, 
    85.49708, 78.09265, 78.93178, 80.02951, 75.44234, 77.29295, 83.8967, 
    86.03164, 84.2664, 91.64489, 94.202, 95.5099, 96.25755,
  98.07093, 98.45152, 98.28407, 97.12589, 96.10219, 95.66692, 95.66119, 
    96.35652, 92.93914, 93.59031, 95.07183, 92.59437, 92.71499, 95.53392, 
    96.91359, 88.32198, 95.01951, 92.53731, 91.10414, 93.01703,
  98.14947, 98.39157, 98.08472, 97.76112, 97.74094, 97.80897, 96.82726, 
    96.15847, 94.24159, 95.31444, 96.38295, 97.57929, 98.28519, 98.10843, 
    97.76981, 97.96198, 98.46796, 98.98096, 98.87282, 99.26506,
  97.52412, 97.65865, 97.57233, 97.63602, 97.55106, 96.88342, 95.80647, 
    94.83234, 94.89419, 95.50294, 96.31863, 96.59122, 96.43008, 95.71189, 
    95.2207, 95.35873, 95.01518, 95.21815, 95.26439, 94.94003,
  96.38762, 96.41242, 96.37945, 96.03471, 95.48445, 94.68688, 93.93958, 
    93.26933, 93.27715, 93.51486, 93.67255, 93.92436, 94.23588, 94.40439, 
    94.21439, 93.42767, 91.7801, 90.8398, 90.92984, 91.1269,
  94.04073, 93.24048, 92.67847, 91.99808, 91.21053, 89.27639, 85.38556, 
    80.93745, 76.82658, 73.98858, 71.44336, 69.96269, 70.43283, 72.74342, 
    75.22315, 76.90775, 78.74753, 81.84843, 83.55633, 82.33005,
  84.63268, 83.21587, 81.37424, 79.36075, 76.96252, 73.86524, 70.05539, 
    68.11713, 67.4997, 67.18499, 66.67027, 66.55957, 67.19302, 68.48689, 
    70.4258, 72.22503, 72.8037, 73.18377, 73.71695, 72.43939,
  79.44804, 78.5481, 77.14573, 75.43469, 73.71008, 71.89384, 70.58235, 
    70.51521, 71.09776, 71.95548, 71.8303, 71.77716, 72.3069, 73.37986, 
    74.70596, 75.70228, 75.40595, 75.55185, 76.11875, 76.53401,
  80.60712, 79.88531, 78.45854, 76.79303, 73.18001, 69.68457, 67.89635, 
    68.08083, 68.86708, 70.25181, 71.12859, 72.0401, 73.36096, 74.53315, 
    75.17937, 76.04025, 76.42283, 76.52528, 76.84055, 77.98895,
  80.15244, 79.53838, 76.86746, 72.68317, 68.23212, 66.03178, 65.88033, 
    66.49667, 67.49338, 69.09083, 71.39192, 73.85759, 75.85949, 77.75086, 
    79.35741, 79.8505, 78.18282, 75.58493, 74.83471, 75.60993,
  74.36211, 71.73727, 67.49914, 64.20137, 63.50114, 64.42229, 65.61012, 
    66.8768, 67.35301, 68.45168, 70.98378, 73.71294, 75.62741, 77.15279, 
    78.22022, 77.66406, 74.49896, 71.10476, 68.50141, 67.38261,
  66.91553, 64.39419, 64.41226, 64.89337, 66.4574, 68.9466, 70.08437, 
    67.02732, 62.85294, 61.13189, 61.68768, 64.00903, 66.69405, 68.55771, 
    70.35822, 70.57929, 67.14069, 61.80915, 58.21979, 57.35752,
  70.17818, 71.50507, 71.32067, 71.50221, 71.78527, 69.81954, 65.36829, 
    61.39937, 59.40092, 56.70063, 55.81086, 56.79948, 58.70354, 59.90591, 
    60.76174, 60.39243, 58.43756, 55.80492, 54.45744, 54.82015,
  71.71985, 70.88663, 69.48805, 68.26005, 66.42757, 64.07585, 63.44176, 
    66.57388, 68.18755, 65.63442, 59.6519, 59.51598, 64.31339, 66.31053, 
    65.37313, 63.69061, 62.17116, 60.40152, 60.02581, 60.19965,
  88.9233, 89.23087, 89.84731, 90.30988, 90.8175, 91.28753, 91.93388, 
    92.24829, 90.78333, 91.3142, 91.61966, 91.77058, 92.0621, 92.30032, 
    92.48692, 92.59611, 91.82511, 91.93027, 92.18619, 92.47505,
  84.10778, 85.34937, 86.79195, 88.23061, 89.7559, 91.14815, 92.4255, 
    93.33933, 89.57632, 90.22038, 90.9486, 92.01376, 92.70656, 93.3249, 
    93.87218, 94.26466, 92.9935, 93.89802, 94.37499, 95.1173,
  85.42161, 87.33116, 89.20392, 91.04562, 92.60396, 93.85902, 94.67657, 
    95.15863, 90.35546, 90.97239, 91.27027, 92.27349, 93.34824, 94.17515, 
    95.21815, 95.73302, 95.27756, 96.26811, 97.37438, 98.41045,
  84.45774, 87.02694, 89.54955, 91.53416, 92.95119, 93.75079, 94.36517, 
    94.56355, 92.41085, 93.41533, 95.27113, 96.61852, 97.48115, 98.04567, 
    98.37428, 98.43522, 98.48173, 98.51429, 98.79575, 98.8846,
  80.33272, 83.14782, 85.41669, 86.62053, 87.28954, 87.47001, 86.85261, 
    86.70374, 86.69976, 87.90469, 90.21524, 92.85449, 94.87439, 96.47815, 
    97.89107, 98.70645, 99.84849, 99.92052, 99.85908, 99.49205,
  79.77958, 80.97922, 81.27213, 81.2765, 81.72195, 82.87323, 84.18768, 
    85.18649, 81.62466, 82.92704, 84.24165, 85.67793, 87.10581, 88.834, 
    90.70812, 92.41608, 98.61278, 99.00607, 98.96152, 98.56818,
  94.86532, 92.1479, 90.38705, 88.95042, 88.69658, 89.20798, 89.081, 
    89.15753, 81.69027, 82.8873, 84.23235, 74.5111, 76.11471, 84.85054, 
    86.0733, 83.27805, 92.16075, 95.39272, 97.20972, 97.90646,
  98.40929, 98.3112, 98.03526, 96.62092, 96.94119, 97.74091, 98.18831, 
    98.45824, 95.05437, 95.13672, 96.15575, 93.7491, 94.34451, 97.46754, 
    98.67927, 90.50488, 97.49895, 95.01603, 92.57429, 93.34329,
  97.48009, 97.91686, 97.86777, 97.43051, 96.95112, 96.53085, 96.92304, 
    97.19659, 95.26439, 95.47592, 96.00858, 96.61341, 97.17518, 97.56276, 
    97.45055, 97.55901, 97.27068, 98.54966, 99.20356, 99.28963,
  97.12584, 97.32555, 97.24536, 97.06476, 97.01997, 96.68253, 96.16327, 
    95.98625, 95.2985, 95.52738, 95.68411, 95.6104, 96.07053, 96.11803, 
    95.92828, 95.79211, 95.88792, 96.15064, 96.58187, 96.61571,
  96.06177, 96.14051, 95.92835, 95.68529, 95.39424, 94.90096, 94.69756, 
    94.99626, 95.00108, 95.07426, 95.15918, 94.75218, 94.41676, 94.29408, 
    94.24331, 94.16579, 93.30569, 93.00463, 92.15999, 91.37746,
  94.64019, 94.2486, 93.51656, 92.33252, 91.71679, 92.33671, 91.34754, 
    89.82322, 88.12925, 86.58539, 84.38276, 81.8605, 81.01997, 82.45937, 
    85.22758, 88.37309, 88.57197, 88.446, 88.12685, 87.77937,
  89.19395, 86.11874, 83.42239, 81.00095, 79.49541, 77.33024, 74.20924, 
    72.22068, 70.88264, 69.4561, 67.49726, 66.58433, 66.73509, 67.92162, 
    69.53728, 71.00904, 71.93073, 73.09869, 74.07906, 73.96928,
  79.66181, 78.55164, 77.38237, 76.08677, 74.34634, 72.43629, 70.79613, 
    70.35958, 70.36, 70.83803, 70.65687, 70.7238, 71.78663, 73.86504, 
    75.22448, 75.85452, 75.28485, 75.55738, 76.35572, 76.8483,
  82.34767, 81.78085, 80.11475, 77.80868, 73.78928, 69.64867, 67.25536, 
    66.86897, 67.54083, 69.06131, 70.87018, 72.776, 74.90812, 76.54937, 
    77.01009, 76.9884, 76.63387, 77.00727, 77.88333, 79.57528,
  80.9649, 80.41373, 76.79929, 72.33906, 68.0905, 65.41259, 65.08944, 
    66.19486, 67.79668, 69.86414, 72.22755, 74.32219, 76.0479, 77.48547, 
    77.82209, 78.22932, 77.68021, 76.46146, 76.40284, 77.61812,
  72.45595, 70.31238, 66.28056, 63.87208, 63.50016, 64.51012, 66.20777, 
    68.29723, 69.9823, 71.04975, 72.36864, 73.65691, 74.7657, 75.61148, 
    75.73898, 75.66598, 73.8351, 71.66631, 70.10436, 69.3441,
  65.09211, 63.99596, 65.65408, 67.64206, 69.37948, 71.52137, 72.07463, 
    68.93452, 64.74879, 63.07943, 63.57972, 65.2305, 67.22133, 68.37933, 
    69.03371, 68.54008, 65.43977, 61.80434, 59.70919, 59.32654,
  74.42589, 76.95261, 77.69005, 77.67079, 77.54314, 75.19813, 69.47266, 
    64.35135, 61.33688, 57.9741, 56.32015, 56.64139, 58.18785, 59.22025, 
    59.46568, 58.6702, 57.05178, 55.7687, 55.51888, 56.03928,
  80.20561, 80.09399, 78.26134, 75.23889, 73.00003, 70.34473, 67.42813, 
    64.59454, 64.71033, 62.30288, 58.59886, 58.15235, 62.69079, 64.89244, 
    63.98616, 62.82234, 62.06502, 61.85314, 62.19275, 63.02562,
  90.81885, 91.02793, 91.49561, 91.63515, 91.96676, 92.38766, 92.60599, 
    92.94988, 91.48125, 91.77053, 92.18018, 92.41044, 92.66595, 93.08168, 
    93.35544, 93.58963, 92.77683, 92.99953, 93.16655, 93.33858,
  86.88527, 87.68816, 88.55054, 89.4461, 90.3929, 91.24829, 91.97926, 
    92.80853, 89.35015, 90.08958, 90.89814, 91.9398, 92.60184, 93.6014, 
    94.37237, 94.89693, 93.27241, 93.96389, 94.56644, 95.10236,
  82.83324, 84.05167, 85.29465, 86.40418, 87.3811, 88.35831, 89.22387, 
    90.09079, 86.09122, 87.13517, 87.77242, 88.53938, 89.4732, 91.00701, 
    92.4156, 93.90515, 93.32491, 94.52322, 95.42452, 96.13477,
  81.19528, 82.36083, 84.02082, 85.49788, 86.63077, 88.23637, 89.56015, 
    90.73872, 88.54084, 89.88107, 91.54932, 93.21055, 94.44515, 95.35973, 
    96.14958, 96.86488, 97.53042, 97.61957, 97.50946, 97.18615,
  76.2764, 77.34199, 77.39141, 78.77201, 80.9102, 83.01244, 84.77303, 
    85.59721, 84.45165, 85.88943, 86.82116, 88.25797, 90.32195, 92.26773, 
    93.89613, 95.26244, 99.1011, 99.33176, 99.09185, 98.31548,
  75.19356, 76.88212, 78.9275, 80.63322, 82.14268, 82.83342, 82.96085, 
    83.01835, 78.70398, 78.8876, 79.54534, 80.67372, 82.04722, 83.66122, 
    85.48432, 87.303, 95.34532, 96.42973, 96.89407, 96.54912,
  90.02301, 86.86197, 86.24605, 86.17915, 86.52344, 86.4917, 85.94597, 
    84.96799, 77.05425, 78.10191, 78.79076, 71.10574, 72.32008, 79.54769, 
    82.5773, 79.59938, 88.47961, 91.87816, 94.29011, 95.47253,
  95.49678, 95.94534, 95.76694, 94.9981, 95.54772, 95.33415, 95.26243, 
    94.991, 90.60494, 90.86838, 90.70062, 89.78182, 90.16773, 93.50262, 
    95.52474, 83.99129, 93.23514, 90.92091, 89.14268, 91.21519,
  95.1523, 95.17796, 95.03745, 94.77127, 94.62218, 94.06455, 93.3825, 
    92.43337, 90.59991, 91.79647, 92.9138, 93.58958, 93.68401, 93.59098, 
    93.22284, 93.81005, 94.07146, 95.02468, 94.38578, 96.50025,
  95.4183, 95.15, 94.84113, 94.92518, 95.07133, 94.69774, 93.69437, 92.20606, 
    90.86947, 90.64603, 90.94102, 91.85176, 92.34554, 91.91196, 91.84256, 
    92.15731, 93.43179, 94.73373, 95.20329, 95.44476,
  95.00365, 95.09772, 95.06727, 94.90132, 95.00122, 95.05318, 94.79961, 
    94.21313, 93.22009, 93.08048, 92.93549, 92.80626, 91.91652, 90.86726, 
    90.02057, 90.32076, 91.28607, 92.26707, 92.86216, 92.8817,
  94.10207, 94.11038, 93.82305, 93.44644, 93.47972, 93.43834, 93.09429, 
    92.70328, 91.25874, 90.78653, 89.61968, 88.4834, 87.7227, 87.67479, 
    89.03704, 89.13937, 90.0373, 89.94182, 90.21942, 89.75679,
  89.14369, 89.06873, 88.45201, 86.73943, 85.02608, 81.53994, 76.81399, 
    74.13633, 72.56419, 70.36341, 67.31918, 65.69302, 66.17966, 68.81259, 
    72.04641, 73.73322, 74.84399, 75.60338, 76.02739, 75.71183,
  84.16984, 83.13777, 81.49061, 78.55196, 74.7224, 71.41392, 69.52742, 
    68.90469, 68.68604, 68.74027, 68.34059, 68.17966, 69.17601, 71.70445, 
    74.75887, 75.78333, 75.32761, 75.16824, 75.80995, 76.74702,
  85.34373, 84.2051, 81.85078, 78.63059, 73.5678, 69.16537, 66.96423, 
    66.66385, 66.8639, 67.8437, 69.31332, 71.20509, 73.51185, 76.03942, 
    77.57133, 77.6729, 77.01482, 76.83215, 77.90915, 80.7748,
  83.0456, 81.55171, 77.17276, 71.863, 67.51836, 65.32428, 65.01808, 
    65.69953, 66.87587, 69.15867, 72.44441, 75.77789, 78.32473, 80.14777, 
    80.72132, 81.20608, 81.21218, 80.26971, 80.45998, 82.08988,
  77.9884, 74.43596, 69.26869, 65.6319, 65.02943, 65.48132, 66.21098, 
    67.29954, 68.47958, 70.32841, 73.39738, 76.92808, 79.65114, 81.15996, 
    81.48135, 81.51821, 80.6218, 78.44938, 76.35175, 74.99828,
  70.28922, 66.75483, 67.04662, 68.96535, 70.09432, 71.30268, 70.62098, 
    66.68952, 62.31601, 61.154, 62.92572, 66.67662, 70.88792, 72.67032, 
    73.79878, 73.91466, 70.7253, 65.69399, 62.5796, 61.94859,
  69.81908, 71.12827, 71.80407, 72.50539, 72.24607, 70.23277, 65.23185, 
    60.98563, 57.87368, 54.78972, 54.02837, 54.97633, 57.42476, 58.86417, 
    59.86999, 59.94035, 58.80054, 57.64978, 57.9587, 59.48024,
  70.93345, 70.54515, 68.99348, 67.32037, 66.72121, 65.24413, 62.85188, 
    61.8453, 61.2878, 58.91481, 55.67495, 55.4176, 60.18477, 63.97275, 
    65.25087, 65.13424, 64.72609, 64.61925, 66.02686, 68.42,
  89.23094, 89.58243, 89.92407, 90.26631, 90.59372, 90.98895, 91.24435, 
    91.58378, 90.05568, 90.33064, 90.60287, 90.8839, 91.14911, 91.45424, 
    91.75216, 92.04765, 91.26154, 91.51596, 91.75218, 92.00089,
  82.70354, 83.21756, 83.98265, 84.75166, 85.76561, 86.61409, 87.44636, 
    88.231, 84.99738, 85.87823, 86.93146, 87.98531, 88.95831, 89.94726, 
    90.91418, 91.99938, 90.55252, 91.631, 92.50856, 93.35786,
  82.21514, 83.07706, 84.12007, 85.1168, 86.18054, 87.5265, 88.77596, 
    89.99638, 85.97659, 87.28983, 88.44821, 89.67381, 90.74081, 91.99686, 
    93.51404, 95.0949, 93.52535, 94.56057, 95.47212, 96.08598,
  85.27638, 87.03573, 88.31702, 89.08487, 90.20966, 91.94239, 93.32045, 
    94.39967, 92.04914, 93.05943, 93.6953, 94.08074, 94.70277, 95.31611, 
    95.79949, 96.14651, 96.99581, 97.06512, 97.1143, 96.8937,
  83.07619, 84.92146, 86.87404, 88.90764, 90.64178, 91.97607, 92.97084, 
    94.09494, 93.30299, 93.60741, 94.12756, 94.28365, 94.45466, 94.23418, 
    94.36032, 94.43735, 97.97073, 97.81476, 97.51375, 96.97801,
  82.9982, 84.50339, 85.94585, 87.2184, 88.49091, 89.36462, 90.10957, 
    90.73736, 86.69846, 86.66, 86.36433, 86.52203, 87.01662, 88.10258, 
    89.58688, 91.08208, 97.43399, 97.97399, 98.24415, 98.18671,
  88.3243, 86.47848, 86.02382, 86.74895, 86.98141, 86.96127, 86.81348, 
    86.21904, 78.7692, 79.69276, 79.68924, 78.20528, 80.00082, 85.18951, 
    86.96627, 85.50588, 92.79226, 94.7069, 95.84191, 96.0397,
  90.10843, 89.79193, 89.55293, 89.89805, 90.91868, 90.8754, 90.25321, 
    89.18371, 83.78607, 83.02711, 79.61321, 82.9732, 84.59555, 90.28412, 
    90.61905, 79.60651, 90.82623, 93.24416, 92.312, 93.66576,
  95.38413, 94.77191, 93.2778, 92.20161, 92.12796, 92.26228, 92.34276, 
    92.60254, 91.30573, 91.66652, 91.76439, 92.20502, 92.10435, 91.00652, 
    91.60231, 92.72901, 92.62679, 94.59547, 93.87337, 94.50394,
  95.85077, 95.80153, 95.59147, 94.66615, 94.62336, 94.3532, 93.72657, 
    93.34023, 93.3379, 93.58755, 93.1698, 92.91661, 93.15273, 93.37738, 
    93.86902, 94.45051, 94.99275, 95.29554, 95.81673, 95.96223,
  94.85394, 94.8771, 95.12621, 95.13659, 94.86644, 94.93243, 94.87921, 
    94.67596, 94.66622, 94.49477, 93.83781, 92.98689, 92.45569, 92.26823, 
    92.31612, 92.77991, 93.14267, 93.21086, 93.10538, 92.74915,
  93.92933, 94.02209, 94.16274, 94.58833, 94.67436, 94.69843, 94.84908, 
    94.90895, 94.42936, 93.68221, 92.31466, 90.88869, 90.18069, 90.40109, 
    90.53242, 90.7625, 90.93346, 91.17306, 91.15208, 90.58834,
  91.06684, 91.07549, 91.00785, 90.70525, 90.17729, 88.65086, 86.02898, 
    84.42305, 83.32923, 81.00953, 77.66313, 75.75375, 76.68663, 79.86283, 
    82.31117, 83.5031, 84.12298, 84.37916, 84.27207, 83.75533,
  88.75135, 87.97975, 86.70975, 84.37808, 81.2725, 78.88288, 77.97638, 
    78.23801, 78.31136, 78.23364, 77.696, 77.91883, 79.42344, 81.62488, 
    83.44154, 83.83673, 83.3642, 83.63732, 84.87625, 86.2104,
  89.04874, 87.91047, 85.16961, 81.91014, 77.44374, 74.07456, 73.36969, 
    74.37971, 75.44872, 76.90646, 78.65342, 80.8856, 83.59219, 85.78842, 
    86.75961, 86.9369, 86.29745, 85.84837, 86.39527, 87.9447,
  86.14996, 84.73193, 80.32545, 75.56693, 71.96404, 70.85977, 72.05404, 
    74.12347, 75.90866, 78.17605, 81.34206, 84.21725, 86.15015, 87.51686, 
    87.5265, 87.40569, 86.83167, 85.91343, 85.60715, 86.28382,
  80.14358, 77.29956, 73.06087, 70.63332, 70.54341, 72.23057, 74.19547, 
    75.61383, 77.01631, 78.98446, 81.17578, 82.94495, 84.18301, 85.01402, 
    84.62705, 84.23242, 83.10167, 81.29288, 79.44102, 77.99909,
  72.40427, 71.06918, 70.95217, 71.69042, 72.56318, 73.86213, 74.65091, 
    72.25996, 69.62221, 69.07681, 70.04399, 71.85958, 73.42373, 74.02989, 
    74.40338, 74.50337, 72.43877, 68.86533, 66.34334, 65.68639,
  68.02939, 69.92538, 70.65508, 70.81649, 70.695, 69.9622, 66.56465, 
    63.87784, 61.95456, 59.53852, 57.64846, 57.49511, 59.13569, 61.45952, 
    63.7794, 64.46069, 64.04018, 63.42901, 64.13804, 65.53073,
  64.57227, 65.54646, 64.81988, 64.74505, 65.37971, 64.62885, 63.30731, 
    63.40771, 65.19331, 64.42033, 59.83017, 57.99878, 62.35824, 67.14597, 
    68.95817, 68.94567, 69.17648, 70.11317, 71.226, 72.1741,
  91.32683, 91.65236, 92.01086, 92.37616, 92.76907, 93.10252, 93.46062, 
    93.95195, 92.50819, 92.69139, 92.76908, 92.94147, 93.02744, 93.11807, 
    93.19417, 93.25938, 92.32297, 92.45924, 92.32648, 92.52626,
  84.63618, 85.41836, 86.42905, 87.44913, 88.4765, 89.44386, 90.45273, 
    91.47756, 88.04768, 88.84692, 89.46891, 90.04284, 90.62283, 91.2738, 
    91.90578, 92.26112, 90.13091, 90.63748, 90.90301, 91.30578,
  80.13895, 81.16997, 82.4883, 83.7728, 85.00661, 86.43305, 87.45718, 
    88.59346, 84.67778, 85.39667, 86.29845, 87.29053, 88.37111, 89.43076, 
    90.56094, 91.43333, 89.7081, 90.37066, 90.91361, 91.23666,
  81.06906, 82.7284, 84.26765, 85.48261, 86.71619, 87.73576, 88.60529, 
    89.41644, 86.35896, 86.745, 87.00259, 87.31982, 87.62765, 87.75849, 
    87.54359, 87.73769, 88.64788, 88.80832, 88.62563, 88.26591,
  81.82959, 84.27401, 86.12012, 87.73405, 89.1513, 90.67792, 91.46712, 
    92.20488, 90.06712, 90.36908, 90.35503, 90.34579, 90.12453, 90.08253, 
    89.55237, 88.55502, 93.11122, 92.28065, 91.41254, 90.15726,
  82.43964, 84.76509, 86.96037, 88.23929, 88.96128, 89.45151, 89.8504, 
    89.92468, 85.30402, 85.46074, 85.90623, 86.45276, 87.11024, 88.28902, 
    89.04957, 90.05096, 96.61916, 96.52478, 96.09386, 95.18942,
  87.70744, 84.85299, 83.48771, 83.31628, 83.15174, 82.89188, 82.30349, 
    81.19691, 72.97638, 72.08539, 70.99758, 73.03337, 74.81312, 79.62646, 
    80.86544, 83.58495, 91.94539, 94.27727, 95.58743, 95.95663,
  93.1368, 92.88615, 92.43037, 91.6509, 90.86686, 90.01511, 88.83864, 
    86.20573, 76.56347, 73.28576, 71.38519, 78.99149, 82.19511, 88.95419, 
    82.24232, 79.61999, 81.29929, 92.94521, 92.40477, 93.56252,
  93.58811, 92.48045, 91.74969, 91.47788, 91.13279, 90.77898, 90.09498, 
    88.73694, 85.37857, 84.45574, 84.92022, 86.64809, 89.03912, 91.19546, 
    92.59772, 93.4829, 93.69661, 93.46191, 93.31726, 94.83891,
  95.16267, 94.71597, 94.03278, 93.63759, 93.10285, 92.63568, 92.09268, 
    91.42652, 90.71054, 90.0545, 90.00418, 90.89987, 92.24951, 93.73891, 
    94.99264, 96.04711, 97.12811, 97.89925, 98.28795, 98.16601,
  94.8217, 94.86457, 94.91579, 95.05254, 95.35038, 95.42065, 95.2121, 94.683, 
    93.82681, 93.53372, 93.04348, 92.25904, 91.64608, 91.56946, 91.67202, 
    91.88865, 92.96978, 93.81672, 94.39129, 94.58696,
  93.45678, 93.71001, 94.04739, 94.4707, 94.98122, 95.04292, 94.34519, 
    92.91418, 91.7391, 90.68533, 88.78039, 87.80866, 87.14192, 86.73573, 
    86.74415, 87.21306, 89.13738, 90.8491, 91.74897, 91.68391,
  90.38747, 90.29236, 90.27374, 90.22741, 89.37988, 86.93858, 83.9221, 
    82.67477, 83.26289, 83.35735, 81.86806, 81.24878, 82.06243, 83.75288, 
    86.13744, 87.79196, 89.52204, 90.67675, 91.54585, 91.61637,
  90.03925, 88.48363, 86.48259, 82.98188, 78.85791, 75.55386, 73.91796, 
    74.52505, 76.55244, 78.64126, 79.43523, 80.03069, 81.31786, 84.06263, 
    87.18984, 88.9464, 90.15134, 91.25169, 92.29271, 92.95812,
  88.95841, 87.2111, 84.1366, 79.96896, 74.8624, 71.08899, 70.20171, 
    71.85658, 75.22957, 78.51829, 81.2224, 83.82038, 86.65837, 88.89183, 
    90.35789, 91.56662, 92.14397, 92.02332, 92.70239, 93.7859,
  84.20676, 82.42442, 77.73499, 72.96694, 69.58995, 68.87637, 70.54932, 
    73.55013, 76.93784, 80.65957, 84.22052, 87.21312, 89.39941, 91.12326, 
    91.99004, 92.27687, 92.19138, 91.5468, 91.82262, 92.18751,
  77.72434, 74.97119, 70.83316, 67.90902, 68.36823, 70.49376, 72.94382, 
    75.24709, 77.86544, 80.68121, 83.31982, 85.66682, 87.47572, 88.8045, 
    89.11187, 89.0658, 88.34238, 87.24846, 86.58752, 85.62944,
  71.67262, 70.1309, 70.06496, 71.11524, 72.46181, 73.20794, 72.9494, 
    70.62759, 68.06246, 68.30467, 70.45688, 74.19415, 77.96494, 79.93561, 
    80.91445, 81.32379, 80.14793, 78.6009, 77.542, 77.09084,
  69.83915, 70.89999, 71.82904, 72.10657, 71.57928, 69.02913, 64.70878, 
    60.82437, 57.2995, 56.12344, 57.28521, 60.53425, 65.55025, 68.99478, 
    70.42453, 70.71621, 71.62167, 72.16182, 72.98094, 73.31422,
  67.94196, 69.01694, 68.23392, 66.10123, 65.09235, 63.58443, 61.95238, 
    59.60825, 61.03472, 62.6997, 63.75225, 64.52027, 68.0471, 69.86326, 
    70.37244, 71.22441, 72.98853, 73.90867, 73.77497, 73.45213,
  92.25591, 92.56815, 92.69531, 92.83132, 93.14468, 93.37677, 93.59355, 
    93.85223, 92.20412, 92.37075, 92.50528, 92.69593, 92.80904, 92.59918, 
    93.02048, 93.27063, 92.3078, 92.34732, 92.45461, 92.52551,
  87.28693, 87.85561, 88.44083, 89.12231, 89.74223, 90.34984, 91.03238, 
    91.63753, 88.07949, 88.72027, 89.33585, 89.8075, 90.31281, 90.96727, 
    91.40158, 91.95537, 89.99843, 90.33194, 90.75558, 91.20464,
  83.93832, 84.87072, 85.84908, 86.7524, 87.85314, 88.94514, 89.90048, 
    90.77173, 86.57715, 87.71853, 88.71416, 89.53783, 90.45213, 91.18348, 
    91.81284, 92.41726, 90.40609, 90.8963, 91.26838, 91.72951,
  84.14311, 85.65115, 87.05642, 88.36449, 89.52106, 90.44726, 91.13766, 
    91.85316, 89.07641, 89.99899, 90.35815, 90.91827, 91.6311, 92.17042, 
    92.80472, 92.97386, 93.96801, 94.08755, 94.01669, 93.96695,
  83.72521, 85.86549, 87.85078, 89.60342, 90.50684, 91.38109, 91.95619, 
    92.69621, 91.73082, 91.96749, 91.86224, 92.26788, 92.85954, 93.18275, 
    93.50514, 93.51038, 97.56193, 97.31424, 96.71851, 96.02942,
  84.57734, 87.08585, 88.93102, 90.45996, 91.46214, 91.75123, 91.55888, 
    91.01952, 86.33105, 86.46296, 86.88483, 87.76266, 88.96898, 90.46826, 
    91.60223, 92.72128, 98.44795, 98.78329, 98.82655, 98.67129,
  90.39218, 88.27493, 87.72566, 88.37497, 88.31721, 87.43237, 86.14178, 
    84.96896, 77.09383, 76.78049, 76.36274, 78.63641, 80.36868, 85.46046, 
    86.01067, 86.70499, 93.86822, 96.12534, 97.56438, 98.2067,
  93.11649, 92.55556, 90.84506, 88.14556, 84.96026, 80.84439, 76.63849, 
    73.22292, 66.40434, 67.5379, 71.59527, 82.87579, 86.73386, 89.96807, 
    76.66164, 77.40316, 77.97851, 92.64088, 91.81834, 93.54692,
  85.18816, 85.07169, 84.62587, 83.82117, 82.32811, 79.93384, 78.25686, 
    77.21151, 74.11951, 73.95892, 75.19087, 77.9688, 82.47414, 86.72878, 
    90.25464, 92.03929, 92.17142, 91.22128, 94.19421, 97.10273,
  86.91153, 85.65669, 84.31662, 83.45148, 82.31385, 81.50703, 80.51034, 
    79.58013, 78.97686, 78.36391, 78.78156, 80.18056, 82.63921, 85.64788, 
    88.55695, 90.4082, 92.48476, 94.42188, 95.42519, 95.49613,
  88.60811, 86.8868, 85.25838, 84.19022, 83.48221, 82.94939, 82.74364, 
    82.42688, 82.08128, 81.53413, 81.53731, 81.84281, 82.59816, 83.55467, 
    84.58649, 85.44672, 87.29581, 89.36396, 91.33218, 92.4425,
  89.22025, 88.59405, 88.30202, 88.3079, 87.85944, 86.92164, 85.31868, 
    84.30621, 83.89146, 83.99605, 83.21893, 83.02479, 83.60287, 84.5649, 
    85.07744, 85.56125, 87.54819, 90.35235, 93.03371, 94.0586,
  90.2541, 89.92326, 89.65643, 90.1689, 90.11948, 87.81757, 84.44038, 
    82.63908, 82.88643, 82.89996, 82.47397, 82.78938, 84.36141, 86.35391, 
    87.8634, 88.96873, 90.88866, 92.72838, 94.30042, 94.6771,
  90.65819, 89.83146, 88.75546, 86.42533, 82.86311, 79.80732, 78.21616, 
    78.24844, 79.49604, 80.84238, 82.01044, 83.77627, 85.85708, 88.11024, 
    90.08555, 90.77145, 91.59081, 92.66006, 93.5165, 94.07993,
  90.04419, 88.94387, 86.35667, 82.63898, 78.22044, 74.92267, 74.07454, 
    75.10995, 77.55653, 80.21152, 82.634, 85.42747, 88.0285, 89.67776, 
    90.52267, 90.80642, 91.131, 91.31525, 92.05052, 93.20045,
  87.83723, 86.16382, 81.89513, 77.4246, 74.22736, 73.20131, 74.44981, 
    76.78201, 79.7169, 82.49763, 85.01754, 87.10247, 88.74727, 89.86745, 
    89.95658, 89.66936, 89.32296, 89.05766, 89.95145, 90.68773,
  84.50594, 81.75436, 78.23257, 76.09018, 75.58724, 76.58828, 78.08434, 
    79.39225, 80.56859, 81.92187, 83.4562, 84.53923, 85.44968, 86.60778, 
    87.29587, 86.73714, 85.54656, 84.5483, 84.87542, 85.8183,
  80.61205, 79.61212, 80.17961, 80.82773, 80.9756, 80.08192, 78.54444, 
    75.88705, 72.98712, 72.13406, 73.41245, 76.32326, 79.35369, 81.6573, 
    82.87228, 82.87895, 81.57858, 80.13572, 80.59997, 82.48577,
  76.38238, 78.41021, 79.52013, 78.97742, 77.69041, 74.57719, 71.30923, 
    67.08817, 62.66155, 60.68147, 61.11335, 64.07261, 68.94623, 73.39283, 
    75.84655, 76.55289, 76.96238, 77.72388, 79.24113, 80.56414,
  69.97517, 70.72179, 69.50591, 68.43892, 69.07293, 68.65814, 67.73242, 
    63.93005, 63.80375, 63.44942, 63.78707, 65.77627, 71.55121, 76.46796, 
    77.62315, 77.72184, 78.69954, 80.79461, 82.55141, 82.66981,
  89.45821, 89.69935, 90.03916, 90.25236, 90.64901, 91.0435, 91.32536, 
    91.57448, 90.11362, 90.3151, 90.50768, 90.70264, 90.90812, 91.20468, 
    91.3624, 91.42896, 90.88775, 90.81664, 91.17476, 91.17161,
  84.27956, 85.07301, 85.91943, 86.89703, 87.86725, 88.89026, 89.84274, 
    90.73992, 87.4348, 88.32841, 89.17702, 90.02893, 90.81425, 91.74215, 
    92.69076, 93.54829, 91.79901, 92.46222, 93.10749, 93.77648,
  86.19068, 87.55962, 88.89171, 90.34306, 91.75314, 92.9922, 94.16424, 
    95.13122, 90.79254, 91.69966, 92.48226, 93.15612, 93.77941, 94.55466, 
    95.82954, 96.85758, 95.50592, 96.13054, 96.59664, 97.07775,
  86.66272, 87.8599, 89.3357, 90.81336, 92.34653, 93.5542, 94.44454, 
    95.43736, 93.09081, 93.61229, 93.94551, 93.86621, 94.29652, 95.34621, 
    96.40329, 97.23503, 98.1693, 98.24878, 98.21465, 98.10917,
  84.84915, 86.63895, 88.21849, 89.6166, 91.09142, 92.43628, 93.28928, 
    93.6759, 92.22481, 92.35892, 92.60941, 93.22649, 94.15578, 95.05521, 
    95.56053, 95.98936, 98.6954, 98.56186, 98.25667, 97.59707,
  82.07072, 84.04267, 85.68443, 86.85426, 87.42841, 88.09225, 89.13428, 
    89.78426, 85.72884, 86.3618, 87.30173, 88.2661, 89.15379, 90.24094, 
    91.25366, 92.80815, 98.3214, 98.44882, 98.48808, 98.02567,
  89.17079, 87.65591, 87.5739, 87.63599, 86.38383, 85.78275, 85.95676, 
    86.26228, 79.17014, 79.5196, 78.91108, 78.79772, 80.24179, 86.9596, 
    89.03249, 84.72921, 91.49923, 94.70047, 96.95181, 97.78129,
  89.1001, 85.04838, 80.97623, 76.05994, 71.11652, 68.77981, 67.64832, 
    67.36539, 62.38111, 63.8476, 67.99978, 83.40995, 86.98714, 90.48952, 
    87.05084, 88.18681, 90.61283, 91.91816, 87.33563, 87.74444,
  86.924, 86.38437, 85.51672, 83.96719, 81.85641, 80.68775, 80.19772, 
    78.65032, 74.92484, 74.06138, 74.16602, 76.67857, 81.98649, 85.53148, 
    86.96392, 86.67361, 84.89547, 83.15874, 86.99701, 90.09946,
  88.09197, 87.64436, 86.90784, 85.945, 84.58407, 83.05922, 81.04848, 
    79.21709, 77.84755, 76.8302, 76.66042, 77.68676, 80.38428, 83.75687, 
    85.55136, 86.63956, 87.34187, 87.84742, 88.42435, 88.00623,
  90.35143, 89.19448, 87.85748, 87.0219, 86.36892, 85.36725, 84.69238, 
    83.49236, 82.61122, 81.67717, 81.15514, 81.42682, 82.57496, 84.62778, 
    86.29613, 86.82616, 87.27523, 87.3135, 88.0637, 88.81284,
  91.80508, 91.43228, 90.80696, 90.53065, 90.12117, 89.50505, 89.33193, 
    89.3466, 88.23387, 86.11026, 84.09737, 83.77651, 84.47374, 85.79079, 
    87.00065, 87.18417, 87.68375, 88.5142, 89.63091, 90.34861,
  91.39594, 91.64259, 91.9613, 91.82104, 90.75494, 88.73777, 86.48431, 
    86.38842, 86.57354, 85.47272, 83.7052, 82.80334, 83.09959, 84.65509, 
    86.34454, 87.3489, 88.0723, 88.95538, 89.81722, 89.98743,
  90.66254, 90.03595, 89.53506, 87.52273, 83.96674, 81.31533, 80.49573, 
    81.23227, 81.91498, 82.30574, 82.00022, 82.13552, 83.04755, 84.4368, 
    86.13489, 87.35, 87.40972, 87.50597, 88.65488, 89.64205,
  90.53786, 89.06576, 87.03732, 84.38175, 80.25599, 77.36707, 76.91075, 
    77.88124, 78.98012, 80.3152, 81.9252, 83.42052, 84.50208, 85.04192, 
    85.7878, 86.85166, 87.29082, 87.557, 88.58923, 90.1866,
  88.33783, 86.45097, 82.23842, 78.25243, 75.5103, 75.0816, 76.14691, 
    77.81836, 79.41142, 81.26668, 82.84987, 83.68269, 84.62536, 85.36832, 
    86.29692, 87.19482, 87.84516, 87.62236, 87.97444, 88.28136,
  81.64185, 78.13642, 75.3402, 74.74239, 75.12533, 76.02437, 77.18653, 
    77.9335, 78.04582, 78.5792, 79.4845, 80.83482, 81.94646, 83.10394, 
    84.07223, 84.55233, 84.27753, 82.61308, 81.09738, 81.32761,
  75.66882, 74.42986, 75.44572, 76.10936, 76.64901, 76.35057, 74.28878, 
    70.3882, 66.87429, 66.45328, 68.81525, 72.1617, 75.48026, 77.36893, 
    78.51034, 78.71578, 76.80077, 73.93724, 73.4175, 74.60477,
  75.09648, 76.3505, 77.04373, 76.09458, 74.32676, 71.37421, 67.01711, 
    62.67515, 60.53351, 59.67745, 60.09858, 61.9598, 64.89316, 67.65329, 
    69.47906, 69.4409, 68.52482, 68.20818, 69.35786, 70.45744,
  72.92184, 73.33027, 72.06942, 69.59254, 68.5667, 66.84675, 66.24391, 
    65.00024, 66.74465, 68.50194, 66.6449, 65.1735, 67.17848, 69.85613, 
    70.88251, 70.20544, 69.19581, 69.0795, 69.38925, 69.45075,
  92.67358, 93.09297, 93.45934, 93.8534, 94.35174, 94.70031, 95.08113, 
    95.4071, 94.09109, 94.52349, 94.8521, 94.88998, 95.42259, 95.72473, 
    95.98472, 95.99113, 95.13039, 95.00797, 95.51652, 95.9114,
  88.25665, 89.2653, 90.43034, 91.43321, 92.52844, 93.51183, 94.48135, 
    95.31477, 91.77143, 92.68342, 93.53672, 94.77596, 95.88101, 96.44676, 
    96.84438, 97.12212, 95.36185, 96.01598, 96.5951, 97.04769,
  87.57413, 88.90025, 90.25187, 91.62863, 92.92178, 94.04086, 95.06349, 
    96.04741, 92.10798, 92.85448, 93.56369, 94.0154, 94.36192, 95.16613, 
    96.02519, 96.59889, 95.54227, 96.158, 96.77695, 97.77203,
  84.3399, 86.0088, 87.78232, 89.5573, 91.38966, 93.19479, 94.92313, 
    96.43486, 94.83757, 95.5508, 96.00237, 96.72236, 97.21269, 97.81898, 
    98.57745, 98.89703, 99.14548, 98.99815, 98.81935, 98.80944,
  80.17941, 82.41105, 84.64021, 86.02612, 86.93349, 86.67658, 85.79764, 
    86.13496, 86.51962, 88.86584, 91.20726, 93.2997, 95.36481, 96.30438, 
    96.94302, 96.69004, 98.82119, 98.73512, 98.28211, 97.7777,
  79.04082, 79.922, 81.30795, 82.285, 82.83868, 82.85074, 83.22515, 83.7475, 
    80.177, 81.30034, 82.37634, 83.65166, 84.909, 86.36697, 87.83228, 
    89.32068, 95.56931, 95.81064, 95.26945, 94.18293,
  87.79426, 85.48975, 85.09538, 86.07851, 86.27299, 87.45551, 87.47265, 
    87.98109, 81.72589, 83.41384, 84.35325, 78.33752, 80.0598, 87.5867, 
    91.22746, 88.69722, 94.31583, 95.21169, 95.73161, 95.40437,
  74.06052, 70.47909, 66.88946, 65.03107, 66.40381, 70.06686, 71.62299, 
    75.13441, 72.78113, 76.99519, 82.62043, 84.37943, 87.66208, 92.82705, 
    95.71712, 96.30367, 97.88555, 96.28149, 93.74602, 93.43291,
  73.95673, 69.05124, 64.47708, 60.36441, 58.10449, 57.36696, 57.17902, 
    56.59031, 55.88653, 57.6516, 60.1225, 64.92752, 72.6044, 79.85522, 
    81.60696, 85.26599, 89.22475, 93.63859, 95.35422, 95.50318,
  84.34194, 82.42722, 80.16857, 77.19373, 74.4963, 71.89977, 69.93659, 
    69.11835, 68.92361, 68.9376, 69.61797, 70.83657, 72.57847, 74.55228, 
    76.2159, 77.29037, 78.92414, 80.44709, 82.32014, 83.81506,
  87.86669, 87.09231, 85.66248, 83.74803, 81.71296, 79.82021, 79.00367, 
    78.98822, 79.5733, 80.13097, 80.59734, 80.45766, 80.15123, 80.65839, 
    81.25082, 81.38605, 82.15207, 82.63263, 83.52306, 84.55369,
  88.21258, 88.06777, 87.56055, 86.44737, 85.12935, 84.33328, 83.9707, 
    84.48128, 85.44582, 85.19767, 84.07476, 83.79863, 84.44544, 85.32113, 
    85.93472, 86.02032, 86.66102, 87.35458, 87.86234, 87.14916,
  87.6604, 88.05984, 88.6834, 88.52904, 87.21323, 84.6814, 81.87157, 
    81.32524, 82.24139, 81.83087, 80.99345, 81.27102, 82.69681, 84.89368, 
    87.30577, 88.38238, 88.60597, 88.64557, 88.53077, 87.67612,
  87.324, 86.89251, 86.12849, 83.73483, 79.67726, 76.09473, 74.06132, 
    74.55795, 76.82982, 78.85841, 80.22375, 82.20795, 84.54289, 86.55048, 
    87.80765, 87.82509, 87.09118, 86.94891, 87.81443, 88.37812,
  87.50529, 86.16911, 83.74869, 79.95002, 74.66212, 70.76277, 69.70094, 
    71.39185, 74.70125, 77.96177, 80.66199, 83.48426, 86.13671, 87.16832, 
    87.23216, 87.19882, 86.92661, 86.85614, 88.25523, 89.34672,
  85.3053, 83.55809, 79.03848, 73.87312, 70.44471, 69.6103, 70.82478, 
    73.51787, 77.10175, 80.1134, 82.78854, 85.27176, 86.2319, 85.99098, 
    85.52604, 85.48087, 85.37259, 85.30718, 85.5385, 84.97852,
  78.1458, 75.77005, 72.69238, 71.04472, 71.84257, 73.53628, 75.00065, 
    76.26792, 77.63653, 79.83673, 81.80315, 82.7573, 82.71425, 82.71416, 
    82.76052, 82.2018, 81.2327, 79.96163, 78.65279, 78.39047,
  72.25158, 70.99068, 71.81648, 73.41303, 74.56808, 74.4258, 72.43319, 
    68.19169, 65.01777, 65.37125, 68.06663, 71.03285, 74.09437, 76.27519, 
    77.92324, 77.90834, 75.40939, 72.96509, 72.12586, 73.20088,
  72.93032, 74.23026, 75.01092, 74.78053, 73.72659, 71.97122, 67.88481, 
    62.71117, 60.08783, 58.47296, 58.07029, 59.70335, 64.25085, 68.40534, 
    70.12904, 69.06555, 67.66381, 67.79662, 69.04755, 70.70804,
  69.94642, 70.08809, 69.34856, 68.70675, 69.2841, 69.30873, 68.89995, 
    66.83001, 67.164, 67.26777, 65.02281, 64.19447, 68.27376, 71.33395, 
    71.94978, 70.48944, 69.3211, 70.03338, 71.30484, 71.5823,
  91.87282, 92.57088, 92.95123, 93.33569, 93.56949, 93.90813, 94.44055, 
    94.66683, 93.33835, 93.80898, 94.15006, 94.32932, 94.49274, 94.88821, 
    95.02869, 95.1748, 94.51465, 94.99297, 95.08249, 95.1405,
  83.98273, 85.34669, 86.88397, 88.49069, 90.15336, 91.76699, 93.06731, 
    94.28125, 91.42596, 92.5793, 93.54116, 94.43053, 95.25814, 95.75333, 
    96.42216, 96.96393, 95.8371, 95.92081, 96.21741, 96.79446,
  81.93569, 84.16748, 86.46329, 88.82284, 90.45213, 91.71434, 92.89601, 
    93.48286, 88.83714, 90.0711, 91.24203, 91.8382, 92.31489, 93.1098, 
    94.18282, 94.74722, 93.75942, 94.64175, 95.74073, 96.86001,
  81.52952, 83.99738, 86.70755, 89.37756, 91.62296, 93.49397, 93.876, 
    94.68474, 92.24886, 93.64817, 95.14005, 96.55228, 97.65188, 98.78752, 
    99.31695, 98.69376, 98.14851, 98.06318, 97.97136, 98.10147,
  77.11388, 79.35143, 80.92609, 82.55003, 83.47871, 84.1927, 86.63063, 
    89.78542, 90.67026, 92.43987, 93.37117, 93.57677, 93.86191, 94.56519, 
    95.60863, 96.00442, 98.41814, 98.94016, 99.20002, 99.1913,
  77.18575, 78.66559, 79.87994, 80.98677, 81.64725, 82.40765, 83.84122, 
    85.50414, 82.88669, 84.24526, 85.15565, 86.12647, 86.75435, 87.62325, 
    88.4543, 89.24412, 95.3725, 95.84702, 95.83671, 95.76069,
  87.1583, 85.58852, 85.9837, 87.19021, 88.11114, 89.07751, 89.87412, 
    91.03671, 83.68394, 83.69237, 85.09537, 79.99538, 80.80857, 84.46272, 
    88.6483, 85.86771, 91.75991, 92.57415, 93.12644, 92.51992,
  84.0705, 84.46368, 86.04321, 87.52238, 89.30299, 92.02042, 93.31882, 
    94.16279, 90.08243, 91.23426, 92.71904, 88.68477, 88.13759, 91.02407, 
    95.70294, 94.30312, 96.3212, 95.86671, 96.01738, 96.45573,
  70.34621, 72.03709, 73.42805, 74.35273, 75.08852, 77.45811, 79.60558, 
    79.71198, 77.84823, 79.80051, 81.70056, 85.59482, 89.81814, 92.87519, 
    93.07745, 92.82768, 93.89875, 95.83674, 96.50169, 96.71645,
  73.71641, 72.27953, 70.90213, 68.4939, 66.14084, 64.76465, 64.4435, 
    64.16322, 63.46084, 62.88754, 63.39187, 64.68884, 66.82869, 67.89871, 
    67.12057, 66.6241, 66.94142, 71.31827, 75.8822, 78.55969,
  79.77592, 79.4901, 78.80357, 77.68688, 76.62948, 75.66467, 74.88245, 
    73.99236, 72.68946, 71.6773, 71.13351, 70.55578, 69.96695, 69.42049, 
    68.84003, 68.18415, 67.61405, 67.20837, 67.25286, 68.26254,
  84.09028, 84.43412, 85.05919, 85.10283, 84.64288, 84.13524, 83.35559, 
    82.94254, 81.87699, 80.01378, 77.97267, 77.09673, 77.21751, 77.91729, 
    78.13108, 77.26716, 76.24976, 76.16041, 76.11511, 75.07088,
  88.29815, 88.6996, 89.08468, 89.1648, 88.37238, 86.65403, 84.36361, 
    83.61366, 83.3719, 82.08724, 79.8129, 78.59426, 78.96426, 80.55251, 
    82.34885, 83.06629, 82.16297, 81.4177, 81.06973, 79.82606,
  90.05623, 89.7499, 89.29559, 87.71163, 84.80991, 82.51722, 81.57883, 
    81.88068, 82.25486, 82.54507, 82.3195, 82.49592, 83.48826, 84.88503, 
    85.54852, 85.57816, 83.84768, 82.42843, 82.11864, 82.25189,
  88.89296, 88.55832, 87.18095, 84.84826, 81.30581, 78.93644, 78.79875, 
    80.13445, 81.68703, 82.94083, 84.01906, 85.28551, 86.79442, 87.27767, 
    86.95093, 86.06649, 83.6671, 81.65609, 81.90336, 83.25306,
  84.81181, 84.14401, 81.07776, 77.38639, 75.2782, 75.86366, 78.14512, 
    80.80732, 82.64111, 83.97924, 85.12937, 86.10909, 86.46181, 85.95002, 
    84.50108, 82.99625, 80.88263, 79.43473, 79.8441, 80.59814,
  78.1094, 76.65123, 74.45556, 73.85658, 76.17751, 79.84465, 82.64921, 
    83.91273, 84.14005, 84.75835, 85.03457, 85.10252, 84.50218, 83.41882, 
    81.52872, 79.68387, 76.87991, 74.28391, 73.02994, 73.0228,
  72.37812, 73.66422, 76.60426, 79.50169, 82.08705, 82.97565, 80.64897, 
    74.83722, 70.34868, 69.75864, 71.55755, 74.29639, 76.21713, 75.86786, 
    74.12258, 72.33109, 69.01567, 66.27213, 65.56083, 66.35191,
  74.61221, 77.47781, 78.59961, 78.51448, 77.27602, 74.67554, 69.71441, 
    65.63301, 64.17592, 62.65259, 62.29955, 63.28339, 63.96382, 62.80785, 
    61.35057, 60.206, 60.01298, 61.69196, 63.90517, 65.57204,
  72.9309, 72.53091, 70.43742, 70.3313, 71.60032, 72.17444, 72.93261, 
    71.19881, 72.31768, 71.89018, 67.57666, 64.608, 64.86179, 63.92011, 
    62.31949, 61.76168, 62.93703, 65.02757, 67.01945, 67.97551,
  92.44656, 92.84383, 92.92935, 93.56908, 94.03983, 94.25198, 94.56112, 
    95.29411, 94.23432, 94.66434, 94.90782, 95.36836, 95.81238, 96.08685, 
    96.45193, 96.69649, 95.9167, 96.18075, 96.46008, 96.45879,
  84.03082, 85.61638, 87.26302, 89.09481, 90.80412, 92.43366, 93.71084, 
    94.65791, 90.88329, 91.4413, 92.14693, 93.04758, 93.95517, 94.50805, 
    95.48145, 96.20597, 94.6481, 95.70925, 96.64113, 97.20576,
  79.25873, 82.22514, 85.34636, 88.40155, 90.98497, 92.58775, 93.43802, 
    94.38682, 90.17081, 91.61883, 92.9464, 94.20927, 95.12182, 95.39165, 
    95.71929, 96.00156, 95.53902, 96.30097, 96.9718, 97.48108,
  82.16591, 84.79829, 87.6346, 90.63933, 92.87019, 94.851, 96.10113, 
    96.47225, 93.98399, 93.04236, 92.88811, 93.62553, 95.16169, 96.90612, 
    99.04012, 99.66672, 99.88999, 99.93786, 99.90725, 99.80213,
  79.62002, 81.5111, 83.00574, 83.97919, 84.17301, 84.60802, 85.14496, 
    85.56092, 84.59933, 86.07955, 88.39689, 90.34322, 92.04484, 93.47274, 
    94.01357, 95.43939, 97.67798, 98.16763, 98.56976, 99.07955,
  79.67934, 80.82704, 81.15103, 81.5703, 81.94547, 82.43655, 82.68977, 
    83.77623, 80.97813, 82.48441, 84.14907, 85.45376, 86.7863, 87.86618, 
    88.66776, 90.64222, 96.58455, 98.74387, 99.24017, 98.8568,
  94.32018, 91.57748, 90.62903, 90.70451, 90.45239, 90.37698, 89.83881, 
    88.7206, 80.73638, 82.05426, 84.86704, 75.80985, 77.13371, 85.31324, 
    88.38007, 80.37704, 87.35298, 89.94381, 92.16888, 93.13631,
  96.39644, 95.98512, 96.14034, 95.46065, 95.13084, 95.47371, 95.61009, 
    95.2656, 90.70457, 92.11037, 93.93089, 89.83878, 90.53585, 94.9328, 
    97.49005, 91.83079, 97.03169, 94.01337, 89.11411, 89.37757,
  95.61465, 96.59207, 97.12569, 96.94709, 95.89806, 94.77151, 95.22554, 
    95.60777, 94.25275, 94.43193, 94.52416, 94.47401, 94.08997, 93.58301, 
    92.96394, 93.56726, 95.02016, 97.22041, 97.52137, 96.27156,
  84.94268, 83.27869, 83.66393, 85.28753, 85.99515, 86.5122, 86.63747, 
    86.88831, 88.24027, 89.3474, 89.15266, 90.04335, 91.11146, 91.66034, 
    90.28693, 89.31622, 90.23721, 91.70831, 93.1937, 93.59663,
  73.33475, 72.22015, 71.53971, 71.75264, 71.45044, 69.72922, 70.49509, 
    71.89963, 74.24625, 75.92873, 77.20947, 78.73388, 80.09251, 80.92773, 
    80.82078, 79.95302, 79.11997, 78.88451, 78.24641, 77.0316,
  70.31522, 70.14265, 70.45045, 71.10715, 71.50649, 71.62294, 71.67351, 
    72.51753, 73.94851, 74.32013, 74.76994, 76.49286, 79.39266, 82.17445, 
    83.57037, 83.53389, 83.20221, 83.37407, 82.91099, 80.92443,
  73.02496, 72.68227, 72.63265, 72.98608, 72.74073, 71.75371, 70.62566, 
    71.24397, 73.29344, 74.40112, 74.33475, 74.72702, 76.31953, 79.88393, 
    83.26815, 84.9495, 85.20962, 85.13505, 85.00542, 83.66219,
  71.52133, 71.29674, 71.10885, 70.07081, 67.79384, 65.62489, 64.9796, 
    66.4019, 69.98784, 72.86978, 74.45441, 75.84657, 77.4908, 80.87333, 
    84.35792, 85.77889, 85.49814, 85.18083, 85.08623, 84.8723,
  72.00772, 71.36624, 70.2294, 68.21626, 64.42598, 60.94418, 59.76426, 
    61.65103, 66.0192, 70.53229, 74.11014, 77.02293, 79.98021, 83.14937, 
    85.0609, 85.31197, 84.21116, 82.96208, 83.06352, 84.11002,
  69.82278, 68.13793, 64.55675, 60.02925, 56.60118, 55.68674, 57.29924, 
    61.29748, 67.45415, 73.46394, 77.52058, 80.7833, 83.58862, 85.62457, 
    86.02119, 85.77967, 84.52765, 83.32072, 83.71902, 84.4087,
  62.12898, 58.52252, 54.94336, 53.42435, 54.66825, 58.51208, 63.67033, 
    68.9731, 73.77638, 77.53967, 80.48646, 83.364, 84.99937, 85.93665, 
    86.29482, 86.39003, 85.50716, 84.0279, 82.57275, 81.97508,
  55.82908, 55.0365, 56.56697, 59.77597, 64.0563, 68.05712, 68.47386, 
    65.01095, 63.12319, 64.79552, 69.20635, 74.4315, 78.8215, 81.61958, 
    83.51452, 84.64111, 83.84348, 81.93309, 80.26648, 78.89342,
  57.19108, 59.84109, 63.05433, 65.19146, 65.44312, 62.95398, 60.19689, 
    58.95498, 60.5333, 59.99411, 61.29663, 65.96883, 71.68886, 75.37668, 
    76.55904, 77.23755, 77.94086, 77.70618, 76.49976, 75.23252,
  57.6536, 58.71726, 59.55197, 60.73362, 61.54508, 62.35223, 64.29475, 
    66.21095, 68.22012, 67.89538, 64.85433, 67.21227, 74.86349, 80.1555, 
    79.29488, 78.87921, 79.20602, 78.35213, 76.84334, 74.5486,
  92.79842, 93.15134, 93.55746, 94.00559, 94.5023, 94.75343, 95.02254, 
    95.29887, 93.73536, 94.03098, 94.35494, 94.7052, 94.99459, 95.32655, 
    95.86188, 96.292, 95.78344, 96.11829, 96.43954, 96.50126,
  86.30473, 87.12184, 88.43143, 89.74675, 90.92599, 91.63798, 92.83213, 
    94.089, 90.43527, 91.30727, 91.95412, 92.52409, 93.22477, 93.93126, 
    94.32209, 95.03654, 94.19438, 95.24953, 96.90007, 98.04579,
  87.72511, 89.53418, 91.12212, 92.54795, 93.9505, 94.65145, 95.32741, 
    96.16731, 93.08616, 95.23471, 96.28221, 95.67464, 95.19372, 96.5634, 
    96.85709, 97.45579, 97.76557, 99.15275, 99.87193, 99.95922,
  82.94272, 84.99673, 87.45493, 89.88419, 92.05394, 93.75295, 94.9962, 
    96.69832, 96.26399, 97.72395, 97.98766, 97.11456, 97.48441, 99.79073, 
    100, 99.84052, 99.58719, 99.26463, 98.90611, 98.53787,
  79.28403, 81.84856, 84.52652, 86.88155, 88.94463, 90.74746, 91.78051, 
    92.43365, 91.62139, 91.93861, 91.52282, 89.35915, 88.07139, 89.43424, 
    92.12418, 94.90498, 98.77306, 99.70976, 99.23521, 98.35522,
  81.13773, 82.51054, 83.85865, 85.4311, 86.41823, 86.42443, 86.06089, 
    84.9753, 78.49653, 76.34322, 75.73664, 77.57491, 80.02071, 82.94692, 
    85.87984, 89.20016, 96.9617, 98.33239, 99.11568, 99.15931,
  94.72029, 92.49078, 91.86036, 91.77001, 91.12823, 90.53586, 89.68392, 
    88.916, 79.14025, 78.50425, 79.76929, 69.50886, 71.47341, 81.10169, 
    86.74532, 79.4874, 88.29388, 91.55123, 93.43941, 94.15499,
  99.17863, 97.45831, 96.52055, 96.15373, 96.48038, 96.77055, 96.92843, 
    96.93664, 91.94826, 92.60313, 94.6984, 89.43819, 90.20952, 95.8502, 
    97.31089, 88.72229, 94.95581, 96.59052, 90.02075, 90.8973,
  99.27505, 99.39117, 99.33728, 99.4359, 99.47022, 99.28934, 98.58945, 
    97.9249, 96.07753, 95.69704, 96.32586, 97.87025, 98.45347, 98.56918, 
    98.38605, 98.01785, 98.27052, 98.91929, 98.6396, 97.71685,
  97.80908, 97.80582, 97.64028, 97.73225, 98.06308, 97.76538, 97.6487, 
    97.23111, 97.1341, 97.03905, 97.13663, 97.04474, 96.69448, 96.647, 
    97.06175, 97.35126, 96.96777, 97.34264, 97.98505, 98.29709,
  96.43262, 96.56985, 95.80476, 95.32582, 94.72878, 92.82246, 90.45534, 
    90.28217, 90.22375, 88.95314, 87.78294, 87.37578, 86.91698, 87.48753, 
    88.60937, 86.95879, 83.35891, 80.81061, 80.07033, 80.33461,
  84.26253, 84.0031, 82.88982, 81.41425, 79.21199, 76.41457, 74.20676, 
    73.60886, 73.42068, 71.98468, 70.00988, 69.20721, 69.85676, 71.76165, 
    73.25419, 73.20336, 71.9843, 71.2705, 70.31787, 68.50613,
  84.35754, 83.73213, 82.88776, 82.10542, 80.99909, 79.07632, 76.56655, 
    75.93701, 76.31754, 75.36742, 73.50362, 72.09549, 71.51194, 72.31837, 
    74.47118, 76.04472, 76.27933, 75.96305, 75.24438, 73.91404,
  86.73492, 85.71422, 83.92571, 81.16271, 78.19366, 75.76353, 74.34498, 
    74.32367, 75.52329, 76.89545, 77.54325, 78.40746, 79.32398, 80.61052, 
    82.70103, 83.39768, 82.19178, 81.2955, 81.06276, 80.8819,
  85.23147, 84.26279, 82.0975, 79.0102, 74.59992, 71.00044, 69.4557, 
    70.01218, 72.13518, 75.00167, 77.90082, 81.12272, 83.81018, 85.92693, 
    87.12821, 86.91898, 85.07334, 83.45071, 83.15218, 83.97134,
  83.33202, 82.57661, 78.95776, 73.39284, 68.19356, 65.69982, 65.79927, 
    67.72521, 71.63799, 76.81403, 81.5162, 84.62463, 87.05891, 88.9665, 
    88.81123, 87.32789, 84.39407, 81.59607, 81.2849, 82.01019,
  76.15668, 73.38766, 69.02692, 65.90622, 65.29515, 66.42115, 69.02106, 
    72.73534, 77.18013, 81.2965, 84.37954, 86.54208, 87.90853, 88.40669, 
    87.01513, 84.32645, 80.46729, 76.85564, 74.60572, 73.47912,
  65.90761, 65.44942, 67.85048, 70.27636, 73.0106, 75.40343, 74.47472, 
    69.78394, 66.2461, 66.06007, 68.15757, 72.03629, 75.72952, 77.36052, 
    76.39941, 74.06931, 69.29244, 65.35357, 63.69417, 63.51968,
  66.85123, 69.91314, 73.11236, 74.03619, 72.62743, 67.72728, 63.01038, 
    60.56459, 60.02895, 57.39083, 56.13984, 56.82768, 58.80537, 60.37854, 
    60.87555, 60.98269, 60.82234, 61.00514, 62.04533, 63.17088,
  68.07682, 69.20073, 68.83746, 67.57604, 65.31989, 63.17283, 63.4488, 
    65.95879, 66.20222, 62.58332, 56.44674, 55.3648, 58.49375, 61.96209, 
    63.67943, 64.72853, 66.19879, 67.98995, 69.66801, 70.37135,
  94.02871, 94.39644, 94.8886, 95.34621, 95.70077, 95.87379, 96.0769, 
    96.29447, 95.24384, 95.48237, 95.61806, 95.78499, 96.09949, 96.2576, 
    96.52861, 96.74847, 96.19703, 96.34147, 96.42101, 96.50052,
  87.61619, 89.22185, 90.91911, 92.43639, 93.95042, 95.10201, 96.05202, 
    96.77892, 93.40735, 93.8335, 94.54428, 95.36333, 95.88791, 95.97322, 
    96.4892, 97.19943, 95.73336, 96.84809, 97.39291, 98.15863,
  86.04342, 88.6455, 91.03461, 92.9528, 94.29918, 95.20854, 96.18478, 
    96.67053, 92.49941, 93.20785, 94.51312, 95.46474, 96.8072, 98.04171, 
    98.55745, 98.94925, 98.50862, 98.93812, 99.29699, 99.63381,
  85.20052, 87.85453, 90.34545, 92.14363, 93.42805, 94.50616, 95.47129, 
    96.22791, 94.20956, 95.18456, 96.42555, 97.44717, 98.44379, 99.07539, 
    99.57577, 99.94679, 100, 100, 100, 99.97723,
  81.48707, 83.93046, 85.67535, 87.2556, 88.7175, 91.10564, 92.76528, 
    93.40714, 93.05801, 93.03438, 92.21814, 92.23077, 93.14381, 94.3936, 
    96.29257, 97.59759, 99.18193, 99.45351, 99.46794, 99.47631,
  81.85952, 82.40559, 84.43289, 86.29057, 87.04506, 87.85825, 88.8364, 
    89.26289, 84.47623, 84.01235, 83.61494, 83.99903, 85.85115, 88.13668, 
    90.21721, 92.48789, 97.78391, 98.8467, 99.12975, 98.97288,
  96.59248, 92.27901, 90.85445, 89.86256, 89.66241, 89.35086, 88.6687, 
    87.7299, 79.08868, 79.21774, 80.61134, 75.41253, 76.21564, 82.00201, 
    85.32627, 80.42859, 88.94895, 92.29117, 94.46835, 95.59502,
  98.89567, 98.73129, 98.50029, 97.41766, 97.1265, 97.17155, 97.22741, 
    97.31728, 93.66312, 93.89847, 94.03094, 91.04869, 90.47993, 93.3662, 
    96.24879, 86.01424, 92.704, 92.33261, 88.66898, 90.57361,
  92.58916, 94.178, 94.9966, 95.67138, 95.52951, 94.77116, 94.39275, 
    94.50057, 93.9473, 95.4193, 96.47412, 96.87438, 96.59953, 95.85963, 
    95.57514, 95.98414, 95.55477, 97.05061, 97.52941, 97.95584,
  93.98573, 92.0097, 90.67915, 90.49745, 90.94974, 90.73359, 89.77863, 
    89.39587, 88.98646, 91.98935, 95.37959, 97.12874, 97.41816, 96.51034, 
    96.06982, 96.13951, 95.7575, 95.94065, 96.35296, 97.03313,
  95.32146, 95.66722, 95.27881, 95.33933, 95.77569, 96.13972, 95.94247, 
    95.25004, 94.13527, 94.00498, 93.23151, 92.57353, 92.82923, 93.94241, 
    93.95988, 93.98456, 93.53805, 93.09261, 93.04723, 92.91223,
  92.22061, 92.90851, 93.0076, 92.08356, 91.83999, 89.25361, 84.76707, 
    81.06448, 76.06073, 67.97938, 63.8992, 62.36841, 64.33131, 68.6123, 
    73.63982, 78.51142, 81.5351, 83.51987, 83.69512, 80.91402,
  71.70894, 71.72581, 69.82426, 68.51373, 65.81334, 62.56011, 58.86984, 
    57.29683, 57.72655, 57.95295, 58.23859, 59.44578, 61.7238, 65.12492, 
    69.53716, 72.79459, 74.54752, 75.1897, 74.88502, 72.98524,
  72.49102, 71.6418, 70.33571, 67.98505, 65.00617, 62.56684, 60.9335, 
    60.79099, 62.08069, 63.75458, 64.88899, 66.16646, 67.99642, 70.24072, 
    73.17151, 75.45107, 76.11353, 76.36433, 76.77349, 77.12105,
  76.8642, 76.39503, 74.75961, 71.88071, 67.35791, 62.99802, 60.64558, 
    61.15114, 63.33887, 65.52424, 67.29488, 69.21875, 71.37888, 73.20406, 
    75.13312, 76.80742, 77.43073, 77.00492, 77.50637, 79.70607,
  78.04131, 76.94001, 73.1371, 67.04928, 61.0746, 57.90893, 57.65697, 
    59.75623, 63.54542, 67.54976, 71.43624, 74.44466, 76.48949, 78.63826, 
    80.34447, 80.38047, 79.0362, 77.21426, 77.66509, 79.74433,
  74.16003, 69.76087, 63.88382, 59.45677, 58.29483, 59.1012, 61.1185, 
    64.20973, 67.93231, 71.36444, 74.4089, 77.0067, 79.10361, 80.8178, 
    81.13078, 80.11426, 78.25912, 76.29602, 75.04154, 74.72451,
  66.43896, 64.31413, 65.41968, 67.68072, 70.26437, 72.41849, 71.92066, 
    67.97488, 64.35541, 62.35467, 63.1172, 66.63592, 71.31074, 74.51909, 
    75.85886, 75.88207, 73.75989, 70.74709, 68.83752, 68.4224,
  69.6322, 72.59496, 75.61308, 76.52343, 75.20762, 69.83036, 63.61406, 
    60.95884, 60.1011, 56.62561, 54.74234, 55.36937, 58.85152, 63.12856, 
    66.01261, 67.40797, 67.18301, 66.34075, 66.33484, 66.65836,
  69.61446, 70.62344, 70.36846, 68.8279, 65.65379, 62.42903, 62.01625, 
    65.70608, 66.39788, 63.50385, 57.17024, 56.78712, 63.64418, 70.11013, 
    72.1094, 72.08168, 71.90567, 71.38019, 71.31575, 70.85493,
  91.6535, 92.02981, 92.45979, 92.83302, 93.29766, 93.59097, 93.87331, 
    94.20892, 93.09088, 93.35371, 93.68668, 94.00538, 94.25137, 94.30057, 
    94.54942, 94.70578, 94.12822, 94.21518, 94.38984, 94.45795,
  85.89604, 87.28609, 88.62013, 89.86685, 91.10684, 92.3103, 93.1535, 
    93.67812, 89.98071, 90.6428, 91.21985, 92.03574, 92.92349, 93.98988, 
    94.78074, 95.39047, 93.71692, 94.03468, 94.56743, 95.41698,
  84.48856, 86.51314, 88.52789, 90.2898, 91.99118, 93.7286, 94.87111, 
    95.12196, 90.0998, 89.58408, 90.09903, 90.20982, 90.33473, 91.41108, 
    91.99017, 92.72337, 92.44808, 93.68594, 95.09057, 96.40454,
  85.27149, 87.75581, 90.03619, 91.93275, 92.72402, 93.78418, 93.99699, 
    93.19676, 90.27837, 91.73022, 93.30913, 94.62373, 95.97409, 97.34208, 
    98.64189, 98.99528, 99.08747, 98.49913, 98.09625, 97.84458,
  81.23847, 83.32778, 84.71249, 82.6175, 80.74292, 81.1771, 82.09495, 
    82.85267, 82.26574, 83.74915, 84.96799, 86.27167, 88.9541, 91.52815, 
    94.00414, 95.7234, 98.76369, 99.5292, 99.23461, 98.82915,
  76.29908, 76.98792, 77.64042, 76.98798, 77.35435, 77.76631, 79.00926, 
    79.75253, 76.46949, 77.39059, 78.33899, 80.1215, 82.35747, 84.69476, 
    87.17987, 89.52943, 96.94878, 98.06203, 98.53814, 98.16772,
  94.35772, 86.73129, 86.31786, 84.74921, 83.15557, 82.12059, 81.55058, 
    82.04832, 75.6431, 77.3295, 77.6097, 69.3575, 72.33872, 81.66996, 
    84.85795, 80.40071, 88.49717, 91.48703, 93.19384, 93.45047,
  98.71098, 98.01536, 97.1414, 95.89048, 96.05759, 95.95933, 96.41673, 
    97.37271, 94.96814, 95.89131, 95.1768, 93.70481, 94.56348, 97.60045, 
    99.34903, 88.22021, 90.71442, 91.30238, 88.71052, 89.27614,
  97.71397, 97.38757, 97.26871, 97.6787, 97.58916, 97.20097, 96.62238, 
    96.12464, 95.04197, 96.08427, 96.92772, 97.94234, 98.48886, 98.69405, 
    99.00479, 99.24812, 98.63674, 99.29126, 97.66825, 98.5532,
  96.50916, 96.68262, 97.24621, 97.71059, 97.60545, 97.23287, 96.87017, 
    96.69579, 96.47768, 94.8995, 94.35587, 94.82531, 95.36417, 95.36434, 
    95.77905, 97.33737, 98.16307, 98.8016, 98.43985, 97.62703,
  96.70415, 96.87048, 97.21602, 97.24815, 97.45346, 97.66085, 97.37927, 
    97.30793, 97.245, 96.45486, 96.00596, 94.84074, 94.51073, 94.09642, 
    94.20853, 94.67049, 94.19141, 94.35796, 93.70855, 92.21321,
  95.52276, 95.59169, 95.45174, 95.6772, 95.67174, 95.6211, 95.17093, 
    94.49499, 93.7822, 88.6826, 81.00192, 75.01267, 73.9357, 78.90614, 
    87.59292, 91.97023, 91.71373, 91.01951, 90.56014, 89.45591,
  90.76508, 90.29018, 88.80994, 86.86868, 84.2183, 78.75761, 71.68559, 
    67.91442, 66.11779, 64.04247, 60.68886, 58.95444, 58.89153, 60.21196, 
    63.45351, 67.20985, 69.29874, 71.04279, 72.24769, 71.95165,
  76.62267, 76.54202, 75.82858, 74.38642, 71.1329, 67.84576, 65.59201, 
    65.18391, 65.73335, 66.58383, 66.44151, 66.11346, 66.57611, 67.99795, 
    69.43843, 70.44775, 70.14175, 70.38924, 70.96861, 71.56583,
  79.10158, 78.58315, 77.11935, 74.77145, 70.57629, 66.63124, 64.42215, 
    64.35695, 65.64512, 67.6446, 69.46474, 71.25603, 72.99838, 74.11526, 
    74.71484, 75.26223, 75.26691, 74.93646, 75.00897, 76.40604,
  79.77505, 79.07152, 76.25671, 71.62975, 66.7403, 63.60803, 62.46926, 
    63.19839, 65.65287, 69.1115, 72.58853, 75.29741, 77.14762, 78.286, 
    79.05887, 79.40042, 78.61819, 77.22791, 77.0288, 78.35244,
  78.4325, 75.18087, 69.69097, 64.84745, 62.87118, 63.10418, 63.85942, 
    65.24564, 67.57949, 69.71477, 71.99982, 74.62685, 76.60078, 78.02663, 
    78.50541, 78.76747, 77.34037, 74.60558, 72.38829, 71.31595,
  69.77689, 66.80733, 66.89091, 68.28965, 69.87635, 71.43913, 71.12874, 
    67.6199, 63.13077, 60.55946, 60.6739, 62.85632, 66.06007, 68.79932, 
    70.88328, 71.77171, 68.92334, 64.65952, 62.00789, 61.11652,
  71.79709, 73.82034, 74.77969, 75.10653, 74.36219, 70.64948, 65.23684, 
    61.49421, 59.22072, 54.5109, 52.21941, 53.05724, 54.81366, 56.1903, 
    57.99546, 59.21944, 59.40079, 59.08091, 59.49375, 60.86945,
  75.2237, 75.77645, 74.80897, 73.02074, 69.57225, 66.62781, 65.11402, 
    65.26977, 66.32326, 61.84004, 55.35796, 54.4719, 58.08511, 60.37209, 
    61.65549, 62.89922, 65.39201, 67.77564, 70.05196, 72.16545,
  91.83558, 92.09624, 92.59961, 92.64895, 93.14893, 93.76616, 94.26466, 
    94.3522, 93.00005, 93.77215, 93.90838, 94.03267, 94.35059, 95.01157, 
    94.8839, 95.22675, 94.39997, 94.58493, 95.02483, 95.25546,
  84.70795, 86.08508, 87.63537, 88.94956, 90.35848, 91.64192, 92.93736, 
    93.9776, 90.64791, 92.16767, 92.71469, 94.08392, 94.2101, 95.39059, 
    95.63911, 96.83201, 95.81814, 96.79051, 97.28311, 98.24215,
  84.41821, 86.23324, 87.33392, 88.89042, 90.4222, 92.5144, 93.72824, 
    94.62561, 89.83714, 91.30247, 92.48664, 94.1808, 95.68591, 97.00462, 
    97.82613, 98.46328, 98.31612, 98.89919, 99.29033, 99.4108,
  83.77001, 85.5893, 87.25066, 87.84945, 88.76477, 90.14706, 91.45995, 
    92.28315, 90.7517, 92.06654, 93.64348, 95.22306, 96.42316, 97.31226, 
    98.08829, 98.51637, 98.97921, 99.05438, 99.07341, 99.02706,
  75.85475, 76.04613, 75.38071, 75.03104, 75.83709, 77.07508, 78.79498, 
    81.32594, 82.88893, 86.10749, 89.18796, 91.31641, 93.51911, 95.47172, 
    96.40242, 96.87101, 99.05491, 99.17404, 99.21983, 99.31653,
  76.07631, 76.13323, 76.87543, 78.44482, 80.07201, 81.31017, 82.05315, 
    82.21758, 78.64142, 79.79121, 81.49216, 83.7018, 85.69601, 87.26535, 
    89.10269, 91.06701, 97.24132, 97.63451, 97.86259, 97.66442,
  93.88212, 90.66388, 89.42058, 88.05078, 87.22271, 87.00863, 86.38396, 
    86.18153, 78.1052, 78.69143, 79.76861, 69.91721, 72.63229, 82.9906, 
    86.85408, 81.39497, 90.17781, 94.09649, 95.9711, 96.9473,
  98.08927, 98.4454, 98.11977, 97.52018, 98.29586, 98.55318, 98.82198, 
    98.74594, 94.62183, 92.59999, 91.65964, 93.32053, 95.29935, 98.64413, 
    99.41053, 84.9012, 92.37208, 93.33426, 87.81148, 89.76144,
  96.1779, 96.69568, 96.73447, 96.57146, 96.65151, 97.18515, 97.18649, 
    96.84631, 95.33148, 95.14846, 95.74123, 96.74361, 97.18343, 97.3179, 
    97.1594, 97.1609, 94.45663, 98.40952, 96.24133, 97.46814,
  95.63847, 95.21732, 95.173, 95.02319, 94.9747, 94.95992, 94.97424, 
    94.88121, 95.0547, 95.49535, 95.69971, 96.39749, 96.57957, 96.68756, 
    96.78685, 96.99928, 96.54151, 96.82735, 97.07002, 97.20325,
  96.21136, 96.60544, 96.61662, 96.6407, 96.80894, 96.86952, 96.8563, 
    96.83844, 96.93366, 96.98679, 96.82924, 96.76752, 96.61474, 96.43179, 
    96.83485, 96.33504, 95.50525, 94.83477, 93.87635, 93.96629,
  94.68696, 94.7478, 94.9496, 95.27943, 95.35517, 95.64198, 95.83704, 
    95.29253, 94.56586, 93.29152, 90.81616, 88.4197, 87.64586, 88.72475, 
    91.15111, 92.05841, 91.92029, 92.03435, 91.66019, 92.32449,
  90.05989, 89.58724, 89.40842, 89.42226, 87.42984, 83.64007, 76.33257, 
    72.44211, 71.39881, 69.90817, 67.25152, 65.6738, 66.20692, 68.4985, 
    71.86319, 75.41192, 77.08827, 78.38743, 80.18954, 81.1599,
  78.30367, 76.90536, 75.17118, 72.55737, 68.87579, 65.5286, 63.15358, 
    62.86394, 64.63467, 66.88329, 67.83473, 68.68073, 70.51473, 73.59743, 
    76.47284, 77.51552, 76.80661, 76.36485, 76.61241, 77.09695,
  80.21078, 79.63094, 77.90506, 74.83362, 70.23034, 65.69574, 63.07454, 
    63.07943, 64.92137, 67.06622, 69.11983, 71.41859, 74.20098, 76.51427, 
    77.62759, 77.78143, 77.57709, 77.47738, 77.87886, 79.49904,
  78.99065, 78.05239, 74.62738, 69.11706, 63.70062, 60.89569, 60.70167, 
    62.32053, 65.28533, 69.38461, 72.95814, 75.90098, 78.11806, 79.2645, 
    79.64101, 80.02445, 79.45881, 77.90173, 77.19804, 78.06818,
  72.0444, 68.63371, 63.45668, 59.12825, 57.63694, 58.75797, 60.68322, 
    62.74677, 65.61856, 69.71805, 73.47751, 76.8712, 79.71504, 81.02464, 
    81.24972, 82.09039, 80.90906, 78.38097, 75.50796, 73.24061,
  60.80304, 58.0998, 57.69441, 58.72909, 61.06782, 64.66357, 66.62623, 
    64.71389, 61.43795, 61.06807, 63.41407, 67.345, 72.19952, 76.26707, 
    78.87157, 79.7364, 76.56957, 71.05537, 66.8826, 64.8371,
  59.97072, 61.88491, 63.13443, 64.73442, 66.17397, 65.32482, 62.18474, 
    59.62305, 57.30681, 54.39269, 54.42231, 57.15672, 61.05021, 65.2085, 
    68.27705, 68.67696, 66.82241, 64.90083, 64.49324, 65.37628,
  63.04803, 63.22806, 63.13544, 62.63471, 60.89418, 59.32324, 59.22252, 
    62.36029, 62.86001, 60.57199, 57.20705, 59.15271, 66.09892, 69.98111, 
    70.71434, 70.34874, 71.03567, 71.94711, 73.53942, 74.65252,
  88.91621, 89.34313, 89.63138, 90.11057, 90.54686, 90.95803, 91.31712, 
    91.65308, 90.42813, 90.77048, 91.15025, 91.51075, 91.91618, 92.08173, 
    92.48446, 92.62699, 91.93118, 92.06757, 92.41496, 92.65768,
  84.69712, 85.80256, 86.90957, 88.00163, 88.9963, 90.01522, 91.05558, 
    92.16019, 89.1133, 90.08347, 91.06859, 92.13449, 93.07356, 93.90977, 
    94.65392, 95.43467, 93.97866, 94.8746, 95.53757, 96.15334,
  83.80042, 85.38614, 86.84308, 88.26103, 89.80602, 91.12984, 92.33656, 
    93.34489, 89.46552, 90.42254, 91.18994, 91.74779, 92.50961, 93.47703, 
    94.57109, 95.64949, 94.69615, 95.47501, 96.23246, 96.86983,
  85.01505, 87.42524, 89.63708, 91.59015, 93.1917, 94.51799, 95.47602, 
    95.98748, 93.56342, 94.23965, 94.90586, 95.19404, 95.64434, 96.23758, 
    96.97675, 97.54491, 98.38222, 98.39834, 98.10406, 97.79068,
  82.90985, 85.6021, 88.40844, 90.24892, 91.6428, 92.80283, 93.7868, 94.6448, 
    93.71742, 94.02428, 94.63785, 95.29676, 96.01017, 96.50788, 96.96245, 
    97.09788, 99.19338, 99.26299, 99.2848, 98.84071,
  81.26371, 84.14009, 86.28887, 87.85565, 88.81373, 89.42573, 90.01025, 
    89.72549, 85.29234, 85.69701, 86.31161, 87.36434, 88.60947, 89.88064, 
    91.36254, 92.67519, 98.14851, 98.30949, 98.19604, 97.41735,
  91.28059, 90.10811, 89.85674, 90.27344, 90.45407, 90.38282, 90.25142, 
    89.20914, 80.73666, 81.25419, 81.77271, 77.64631, 78.8736, 84.20313, 
    86.26677, 84.51356, 91.75452, 94.55952, 95.67236, 96.22743,
  93.73866, 94.96889, 95.50679, 95.41637, 95.47869, 95.42108, 96.18732, 
    95.40812, 90.49742, 90.98736, 89.56306, 87.90565, 88.55003, 92.61905, 
    94.92302, 82.06078, 82.66029, 91.28255, 91.59582, 93.7672,
  96.24654, 95.56821, 94.61498, 94.1829, 93.97156, 93.80475, 93.56828, 
    93.43874, 91.7822, 92.50464, 93.09129, 93.26488, 92.90112, 92.90518, 
    93.29309, 93.96371, 93.93289, 95.64837, 93.68989, 95.03328,
  96.75387, 96.61434, 96.34381, 95.94397, 95.72232, 95.18656, 94.39889, 
    93.2205, 93.37231, 93.57599, 94.1198, 94.19963, 94.31606, 94.88266, 
    95.22849, 95.66335, 96.03126, 96.40943, 96.27946, 96.02554,
  96.49772, 96.61126, 96.66632, 96.64325, 96.60473, 96.40843, 95.83076, 
    94.9249, 94.19458, 94.18443, 94.14793, 94.21188, 94.66112, 94.91972, 
    95.14953, 95.18964, 95.49297, 95.90978, 96.01795, 95.53064,
  95.77234, 95.75259, 95.54315, 95.57235, 95.33785, 94.97838, 94.67425, 
    94.13304, 93.26675, 93.29197, 92.71327, 91.9336, 91.52165, 92.10545, 
    92.28323, 91.80135, 91.53261, 91.56395, 91.88313, 92.01931,
  91.64047, 92.80538, 93.43967, 93.51305, 92.28869, 90.67636, 86.94965, 
    84.42844, 83.15994, 81.39764, 77.94238, 75.08019, 74.80527, 76.11115, 
    77.21626, 78.22938, 78.62339, 78.89857, 79.13703, 78.74298,
  84.22543, 83.51917, 82.38747, 79.62089, 75.09474, 71.2412, 68.91087, 
    68.52881, 68.93747, 69.80541, 69.94329, 70.26092, 70.90737, 72.58791, 
    74.79953, 75.77689, 75.05158, 74.71941, 75.30382, 76.1101,
  82.23995, 81.82243, 80.09113, 77.11543, 72.43379, 68.51073, 66.15771, 
    66.2104, 67.65715, 69.55334, 71.34981, 72.86504, 74.43165, 75.65137, 
    76.32941, 76.50196, 75.66158, 75.38412, 75.78407, 77.56162,
  77.91127, 77.85201, 75.36879, 71.41518, 67.14249, 65.08905, 65.55936, 
    67.63644, 70.1913, 72.84459, 75.4508, 77.11765, 78.21997, 78.48702, 
    78.33942, 78.48777, 77.7007, 76.62155, 76.47974, 77.6538,
  71.82005, 69.97418, 66.198, 63.42335, 63.08128, 64.8606, 67.51638, 
    70.05732, 72.27598, 74.0499, 75.92159, 77.56839, 78.68, 78.8157, 
    78.47062, 78.29227, 77.12856, 75.62635, 73.77906, 71.89193,
  63.85206, 61.89539, 62.28405, 64.44781, 67.11082, 70.12882, 71.9065, 
    70.04185, 66.28038, 64.97694, 65.91505, 67.96777, 70.2286, 71.8139, 
    72.97328, 73.42876, 70.96771, 67.12857, 63.82712, 62.30705,
  65.30927, 66.85506, 67.87708, 70.03157, 71.74117, 70.62167, 66.47262, 
    62.36673, 58.67719, 56.17585, 56.04335, 58.23602, 61.6546, 64.2714, 
    65.67691, 65.76706, 64.03295, 62.01927, 61.35151, 61.8232,
  68.75951, 67.9252, 66.38177, 66.17552, 65.42924, 64.03669, 62.80816, 
    63.56756, 63.47833, 61.8664, 59.35441, 60.45338, 66.72578, 69.83652, 
    70.43968, 69.83991, 69.13391, 68.63446, 68.58353, 68.78962,
  90.39658, 90.69701, 91.03044, 91.37196, 91.74318, 92.08233, 92.40121, 
    92.74551, 91.33734, 91.66987, 92.01801, 92.29074, 92.58064, 92.83862, 
    93.14882, 93.64499, 92.86414, 93.05978, 93.28112, 93.42737,
  83.51214, 84.3993, 85.18129, 86.00459, 86.81953, 87.78151, 88.92296, 
    90.0992, 86.91761, 88.00384, 89.08659, 90.08331, 90.99933, 91.76247, 
    92.69919, 93.55968, 91.80088, 92.54365, 93.2803, 93.84602,
  83.04505, 84.20846, 85.46259, 86.61989, 87.62403, 88.85268, 90.00706, 
    91.38213, 87.3014, 88.57983, 89.72028, 90.63808, 91.99221, 93.15948, 
    94.04514, 95.09953, 93.57687, 94.32811, 94.96684, 95.49917,
  84.74532, 85.96754, 87.56065, 88.95861, 90.40382, 91.86485, 93.04565, 
    94.33382, 91.91895, 92.63139, 93.30678, 93.75958, 94.41747, 95.18584, 
    95.90256, 96.40619, 97.50446, 97.51829, 97.2121, 96.78259,
  82.48874, 84.31881, 87.59357, 89.78691, 91.65481, 92.94941, 93.90749, 
    94.61897, 93.30528, 93.90498, 94.32983, 94.8568, 95.36823, 95.7431, 
    96.0633, 96.18756, 99.31107, 99.0779, 98.28702, 97.55078,
  82.02528, 84.60242, 87.93342, 90.29358, 92.02186, 92.98347, 93.27553, 
    93.27001, 89.10327, 89.25814, 89.33611, 89.90287, 90.7397, 92.00066, 
    93.56191, 94.54156, 99.20775, 99.16507, 98.87708, 98.38669,
  91.4769, 89.89333, 89.80304, 90.98008, 91.87702, 92.21752, 91.94707, 
    91.57019, 83.67449, 84.14326, 82.35165, 82.17808, 84.56513, 91.02062, 
    92.38697, 90.67089, 95.96159, 97.20277, 97.95076, 98.39746,
  93.03757, 93.28413, 92.98864, 92.80264, 92.77538, 92.76413, 92.98342, 
    92.97329, 88.72659, 87.6943, 82.70412, 87.20729, 88.69591, 94.26053, 
    92.78545, 82.35762, 86.80605, 95.52929, 95.16953, 96.65072,
  94.69654, 94.16575, 93.82278, 93.85387, 93.66022, 93.56122, 93.32634, 
    93.38426, 91.6172, 91.37441, 91.38244, 91.73931, 91.19955, 90.94865, 
    91.75269, 92.49042, 91.72981, 93.44657, 91.91019, 94.70853,
  96.0211, 95.62247, 95.19515, 95.11488, 94.76974, 94.55254, 94.285, 
    94.43806, 94.34259, 94.77994, 95.2047, 94.78276, 94.23171, 93.68673, 
    93.19209, 93.12495, 92.76086, 92.76011, 93.3056, 93.28261,
  95.54858, 95.20888, 94.87532, 94.95708, 94.94565, 94.8795, 94.77895, 
    94.81919, 94.27075, 94.62815, 95.27145, 95.04939, 94.43222, 93.50324, 
    92.89864, 92.7193, 92.46893, 92.64838, 92.64388, 93.04321,
  94.31447, 93.85197, 93.53511, 93.49442, 93.92883, 94.25967, 94.02968, 
    94.05859, 92.99241, 93.38443, 93.33508, 92.65788, 92.34286, 92.3738, 
    92.37247, 92.40137, 92.46798, 92.58412, 92.1255, 91.8427,
  88.32112, 88.23896, 88.1131, 88.13882, 87.93876, 86.73181, 83.91024, 
    82.99596, 82.36847, 81.53838, 78.90741, 77.21024, 78.19075, 81.49258, 
    84.23248, 85.43086, 85.5566, 86.13219, 86.77297, 86.52804,
  86.86998, 85.89639, 84.59894, 82.11195, 77.80981, 73.78008, 70.72047, 
    69.33756, 69.18495, 70.26067, 70.8617, 71.80652, 73.78236, 77.44662, 
    81.47199, 82.84339, 81.92667, 81.63391, 82.57172, 83.79544,
  84.19284, 83.45213, 81.65516, 78.51546, 73.42305, 68.73705, 65.99162, 
    65.60863, 66.7261, 69.46557, 72.03855, 74.55144, 77.08714, 79.29218, 
    80.93119, 81.5188, 80.79037, 80.51141, 81.73397, 84.49879,
  80.33601, 78.94829, 76.21757, 72.55843, 68.25757, 65.36973, 64.75695, 
    66.35847, 69.1168, 72.43828, 75.75327, 78.71379, 81.09025, 82.95869, 
    83.3454, 83.44179, 83.0787, 82.3502, 82.54863, 84.02607,
  78.76846, 74.99847, 70.55258, 67.36562, 65.92492, 66.14846, 67.36031, 
    68.95325, 70.97925, 73.2662, 75.62144, 78.07415, 80.20487, 81.87356, 
    82.12165, 82.41397, 81.83759, 80.38333, 78.53911, 77.1555,
  76.34728, 71.5443, 69.33578, 69.15428, 70.00188, 71.04212, 71.40874, 
    68.61829, 64.37595, 63.28626, 64.99756, 68.1515, 71.19743, 73.3563, 
    75.05669, 76.18224, 74.27134, 70.71139, 67.98683, 66.63852,
  75.16364, 74.58011, 73.6133, 73.37777, 73.44408, 71.47121, 66.92892, 
    61.80014, 57.22575, 54.33913, 54.51201, 57.45933, 61.39949, 64.96609, 
    67.14708, 67.41098, 65.99292, 64.89837, 65.02725, 65.57329,
  74.03961, 72.7858, 70.84545, 69.84805, 69.12959, 67.06212, 64.57922, 
    61.27417, 60.58335, 58.50672, 56.12529, 58.23113, 64.51389, 68.82112, 
    69.98809, 69.84078, 69.39194, 70.12445, 71.85898, 73.56689,
  92.55531, 92.71696, 92.8677, 93.17818, 93.47694, 93.57288, 93.73112, 
    94.02492, 92.44167, 92.66988, 92.86943, 92.97587, 93.15392, 93.38991, 
    93.4719, 93.54063, 92.67392, 92.85749, 93.20578, 93.3354,
  84.98476, 85.78521, 86.53493, 87.2449, 88.31774, 89.24516, 89.68466, 
    90.22686, 86.73827, 87.53912, 88.29076, 88.98237, 89.64177, 90.58099, 
    91.25618, 92.30971, 90.32104, 90.58266, 91.03526, 91.42345,
  81.77288, 82.59483, 83.68721, 84.39124, 85.10562, 85.87872, 86.76848, 
    87.4166, 83.36212, 84.24009, 85.44041, 86.37716, 87.33311, 88.27388, 
    89.16422, 90.13732, 88.39307, 89.1086, 89.96134, 90.76513,
  82.00342, 83.30904, 84.39165, 84.88066, 85.57037, 85.9133, 86.06606, 
    86.38879, 83.58215, 84.15766, 84.93786, 85.92948, 86.31176, 86.79539, 
    87.02644, 87.51841, 88.73077, 89.22906, 89.43132, 89.29754,
  81.12791, 83.49116, 85.34074, 86.46274, 86.88472, 87.61961, 88.0317, 
    88.94055, 87.84597, 88.06683, 88.52015, 88.97862, 88.881, 89.05303, 
    88.9541, 88.38867, 92.85612, 91.85785, 91.05535, 90.1668,
  81.49863, 84.13483, 86.10122, 87.64706, 88.78649, 89.62411, 90.32277, 
    90.2897, 86.3233, 86.84368, 87.46469, 88.25879, 89.11417, 90.14572, 
    90.94366, 91.6401, 97.42817, 97.07342, 96.57902, 95.83139,
  87.55859, 85.45265, 85.06272, 85.46832, 85.48515, 85.44511, 85.1395, 
    85.25796, 77.47295, 76.38558, 74.67175, 76.88924, 78.68156, 83.00127, 
    84.90247, 87.04731, 94.23872, 96.16063, 96.9964, 97.16771,
  90.75419, 90.86425, 90.98064, 90.92693, 90.34484, 89.78783, 89.04551, 
    87.85944, 79.82394, 76.80342, 73.2382, 79.11162, 81.76905, 88.98428, 
    82.9139, 77.6531, 75.60674, 92.59841, 92.44201, 93.7932,
  94.80997, 93.02282, 91.23315, 89.97105, 89.15179, 88.79929, 88.381, 
    87.44911, 83.00626, 81.33485, 80.29485, 79.49761, 79.4891, 80.88136, 
    83.99838, 86.54047, 86.80999, 84.62563, 88.14315, 91.83263,
  98.04931, 96.0267, 93.19512, 91.07278, 89.94522, 88.51784, 88.28295, 
    88.28497, 88.119, 87.82652, 87.36761, 86.52816, 85.79375, 85.66499, 
    85.91297, 86.77362, 88.34608, 90.5125, 92.34381, 94.03089,
  95.31593, 94.0109, 91.90443, 89.54652, 88.47707, 87.73184, 87.17195, 
    86.85127, 87.25928, 87.53315, 87.93983, 87.66449, 86.51529, 85.72015, 
    85.89988, 87.00023, 88.62294, 90.6433, 92.23841, 93.6041,
  91.35765, 90.47855, 89.69212, 89.05532, 89.32134, 89.33572, 88.1833, 
    86.85391, 86.11488, 86.3504, 86.7915, 86.85526, 86.17325, 85.89874, 
    86.08331, 86.9912, 89.00093, 91.01351, 91.65259, 91.35881,
  91.73537, 91.6625, 91.78303, 92.43797, 92.97321, 92.15279, 89.27561, 
    87.10314, 85.64667, 84.10874, 82.51637, 82.15907, 83.70737, 86.04913, 
    87.11014, 87.09311, 87.822, 88.90046, 89.20612, 88.91866,
  92.58386, 92.831, 92.30756, 90.49129, 87.63802, 85.27254, 83.73443, 
    83.30061, 82.98861, 83.01364, 82.83411, 83.0767, 83.90563, 85.30849, 
    86.92214, 87.20148, 86.40942, 86.6074, 87.72285, 89.1403,
  90.18983, 89.96317, 88.3503, 85.31269, 81.07883, 77.98041, 77.11092, 
    78.27102, 80.4709, 82.58485, 84.02159, 85.34114, 86.26382, 86.63359, 
    86.54277, 86.11004, 85.144, 85.16093, 86.52508, 88.81928,
  84.65511, 84.02796, 81.08858, 77.27917, 73.89108, 72.53003, 73.53649, 
    76.23054, 79.67612, 82.67407, 84.99046, 86.83276, 88.0422, 88.33301, 
    87.40464, 86.62852, 86.01562, 85.43005, 85.57033, 86.37904,
  79.92416, 77.89605, 74.68173, 72.08051, 70.63086, 71.20242, 73.78149, 
    76.2135, 78.33968, 80.1764, 81.95173, 83.66885, 85.31606, 86.19049, 
    85.70641, 84.9874, 83.75769, 82.55784, 81.38558, 80.54636,
  76.69476, 74.78356, 74.29874, 74.1576, 74.43437, 75.65053, 75.92263, 
    73.60139, 70.26009, 69.16545, 71.02705, 74.60734, 78.28608, 80.47694, 
    80.88799, 79.68686, 76.81228, 74.06719, 72.29712, 71.4129,
  76.97889, 78.4296, 78.41375, 77.9688, 77.3409, 75.66761, 71.66557, 67.3802, 
    63.40472, 61.14185, 62.4223, 65.42112, 69.36404, 71.91754, 72.32962, 
    71.17194, 69.55299, 68.75302, 68.42083, 68.4659,
  76.54897, 77.12339, 75.76229, 74.63152, 74.91374, 72.39832, 68.62617, 
    64.40134, 63.95277, 65.02423, 66.55879, 67.67834, 71.32504, 72.69505, 
    71.54419, 70.20616, 69.80437, 70.48985, 71.20747, 71.67169,
  95.03599, 95.35587, 95.65775, 95.90239, 96.14656, 96.33324, 96.54917, 
    96.6296, 95.34806, 95.63989, 95.85228, 95.99699, 96.30082, 96.63667, 
    96.86756, 96.87888, 96.17397, 96.30355, 96.4633, 96.63689,
  90.81054, 91.56707, 92.17435, 92.55547, 93.02737, 93.81364, 94.82986, 
    95.70248, 92.92673, 93.68975, 94.24529, 94.79884, 95.27594, 95.45325, 
    95.68597, 96.07661, 94.13525, 94.51345, 94.9585, 95.35965,
  84.93221, 86.44965, 87.33961, 88.67281, 89.8801, 91.32682, 92.5967, 
    93.65644, 89.6112, 90.37144, 91.30183, 92.08436, 92.79805, 93.20667, 
    93.92612, 95.08137, 93.19981, 93.69128, 94.16975, 94.6348,
  84.0616, 85.85103, 87.20856, 88.73022, 89.90139, 90.98135, 91.85196, 
    92.62065, 90.26391, 91.14333, 91.97487, 92.49596, 93.07107, 93.76991, 
    94.14114, 94.19255, 94.8146, 94.89112, 95.05131, 94.95453,
  84.05151, 86.42181, 88.53938, 90.25166, 91.57564, 92.48091, 93.09828, 
    93.35557, 92.00321, 92.84814, 93.1414, 93.61584, 93.8156, 93.82838, 
    93.77127, 93.94366, 98.02943, 97.95352, 97.76385, 96.68867,
  83.24366, 86.11847, 88.11958, 89.57443, 90.65985, 91.34892, 91.85287, 
    92.08887, 87.78014, 88.03062, 88.43333, 88.92724, 89.59737, 90.51892, 
    91.76947, 92.46136, 98.6568, 98.86671, 98.66122, 97.98404,
  88.03168, 84.71333, 84.41583, 84.94229, 85.02761, 85.03381, 84.79535, 
    84.51179, 76.65884, 75.99855, 75.51528, 76.58595, 77.99998, 82.46215, 
    82.74309, 85.32277, 92.60719, 94.40926, 95.6219, 95.8632,
  89.95269, 88.91312, 87.40188, 85.75729, 84.30712, 83.34695, 82.00143, 
    80.45477, 72.989, 72.24245, 72.27503, 77.12423, 78.96246, 81.6497, 
    71.33067, 74.39124, 76.52115, 92.90733, 93.51434, 95.04353,
  88.77818, 88.25514, 87.76374, 87.35213, 86.44589, 86.34267, 85.86017, 
    84.20986, 80.65682, 80.4155, 81.10086, 81.87988, 83.60418, 85.63268, 
    88.08112, 89.58109, 90.8785, 90.62326, 93.71123, 96.53194,
  87.57196, 85.42584, 83.94308, 83.86304, 84.22832, 84.13718, 83.89201, 
    83.75801, 83.78495, 82.67567, 82.17733, 83.27262, 85.29871, 86.88943, 
    88.10804, 91.40944, 94.40001, 95.72067, 96.41888, 96.41974,
  81.39658, 80.54829, 79.5811, 79.00166, 79.83177, 81.5089, 82.46311, 
    84.56202, 86.1098, 85.19248, 84.27026, 84.5912, 85.43849, 86.34905, 
    87.32876, 88.90539, 91.11465, 92.56589, 93.4773, 93.25801,
  79.69444, 79.03323, 79.32935, 80.62145, 82.25465, 84.24743, 84.9067, 
    85.77876, 86.23248, 86.14083, 85.97594, 86.57257, 87.1609, 87.28873, 
    87.84949, 88.8265, 90.91483, 92.70593, 93.24777, 92.499,
  83.34553, 83.89942, 84.4663, 85.56348, 86.17583, 85.57774, 83.84266, 
    83.49036, 84.69253, 84.45914, 84.02486, 84.96941, 87.05241, 89.03708, 
    90.53841, 91.38076, 91.77147, 92.55989, 93.06865, 92.77996,
  88.00962, 87.82132, 87.03215, 85.00643, 81.16714, 78.0792, 77.1712, 
    78.48001, 81.0463, 82.768, 83.33304, 84.24573, 86.64241, 89.48457, 
    91.77673, 92.20815, 91.2141, 90.93884, 91.89436, 92.92421,
  87.76509, 87.24537, 85.27291, 82.26797, 78.30444, 75.28458, 74.42775, 
    76.00542, 79.20955, 82.03666, 83.74425, 85.53528, 88.12016, 90.68568, 
    92.43133, 92.83488, 91.91535, 91.22578, 91.98408, 93.40396,
  85.68658, 84.60887, 81.79912, 78.67748, 75.96194, 74.86048, 75.41309, 
    77.45581, 80.48763, 83.32239, 85.48281, 87.7571, 90.00603, 91.87565, 
    92.69395, 92.61405, 91.68147, 90.96366, 91.4586, 91.97031,
  82.69319, 80.87682, 78.23476, 76.48805, 75.64062, 75.80701, 77.26395, 
    79.34543, 81.17396, 82.66259, 84.20174, 85.88137, 87.5175, 88.97175, 
    89.19294, 89.02183, 88.17603, 86.90299, 86.42623, 86.03789,
  79.33757, 77.60197, 77.3287, 77.72667, 78.56059, 79.31142, 79.56496, 
    77.6164, 74.19576, 73.28628, 75.21455, 78.07522, 80.71307, 83.02487, 
    84.03724, 84.59192, 83.88129, 82.13966, 81.59652, 81.23518,
  77.68372, 78.70782, 79.71761, 80.39252, 81.00838, 79.5519, 75.30957, 
    69.84837, 66.24357, 63.90884, 64.81832, 68.54417, 74.30099, 77.75349, 
    79.02524, 79.36242, 79.24106, 79.25073, 79.77238, 78.84564,
  75.7466, 76.59883, 76.11191, 75.45445, 74.83285, 72.5173, 69.22556, 
    64.41747, 63.04602, 62.81911, 64.78814, 68.08359, 74.238, 77.51308, 
    77.694, 77.72378, 78.37501, 79.44635, 79.68701, 78.64543,
  93.246, 93.59023, 93.98288, 94.11693, 94.60224, 94.81236, 95.05097, 
    95.59052, 94.05547, 94.47627, 94.72704, 94.87185, 95.37038, 95.14169, 
    95.38651, 95.97153, 95.16191, 94.92908, 95.5163, 95.70068,
  85.98651, 86.92688, 87.85034, 88.79745, 89.9286, 90.91314, 91.97143, 
    92.97105, 89.62832, 90.41274, 91.11901, 91.92464, 92.7906, 93.56302, 
    94.41302, 95.10542, 93.38332, 93.76969, 94.367, 95.02334,
  83.07993, 84.40519, 85.77365, 87.16496, 88.69074, 90.22945, 91.86758, 
    93.11238, 89.17612, 90.42539, 91.47019, 92.507, 93.36706, 94.31192, 
    95.03675, 95.91817, 94.31213, 94.79613, 95.17133, 95.4927,
  83.38744, 85.27511, 86.96353, 88.44036, 89.89676, 91.36097, 92.6692, 
    93.93744, 91.64819, 92.69947, 93.49603, 94.40861, 94.88271, 95.13405, 
    95.52886, 95.94884, 96.74174, 96.61555, 96.05045, 95.48412,
  83.58878, 85.99299, 88.18524, 89.91895, 91.25445, 92.13511, 92.79404, 
    93.26655, 92.239, 92.76459, 93.15497, 93.56695, 93.86913, 94.11043, 
    94.16404, 94.05806, 97.16871, 96.69962, 96.17164, 94.69357,
  83.22335, 85.56571, 87.66842, 89.21179, 90.29386, 91.0071, 91.25975, 
    91.25885, 86.95301, 86.97144, 87.13085, 87.30363, 87.58898, 88.24075, 
    89.13419, 89.74393, 96.69704, 96.82766, 96.56758, 95.50827,
  87.65826, 84.40398, 83.82121, 83.9402, 83.6712, 83.45358, 83.245, 82.93845, 
    75.39621, 74.92, 74.32433, 75.17488, 76.15577, 79.38194, 81.2356, 
    82.22759, 89.83523, 92.18528, 93.48643, 93.67451,
  82.17764, 80.91814, 79.69134, 78.83141, 78.57752, 78.26472, 77.9472, 
    77.14404, 70.23996, 68.2881, 66.23544, 69.12242, 72.39785, 76.43988, 
    71.92876, 74.37578, 80.80209, 87.90955, 88.57774, 90.82788,
  84.5049, 85.79755, 86.88088, 88.09417, 89.29326, 89.78634, 89.19007, 
    87.30301, 82.82898, 81.4498, 80.58875, 80.24088, 81.82577, 85.01622, 
    86.0227, 86.44891, 86.11462, 84.47856, 88.07694, 90.83466,
  80.21158, 82.22968, 84.59439, 86.61396, 87.67709, 87.79792, 87.36675, 
    87.04875, 87.07772, 85.99096, 85.02616, 84.87022, 85.32029, 85.85379, 
    86.3633, 87.51916, 88.97382, 89.98283, 90.27609, 90.21214,
  78.49687, 79.53497, 80.91387, 83.19012, 85.35089, 86.52472, 86.47666, 
    86.46081, 87.3877, 87.49477, 87.44366, 87.54291, 87.75282, 87.90564, 
    87.76188, 87.85262, 88.57665, 89.33745, 89.41021, 88.88509,
  81.11967, 80.141, 80.18185, 81.76521, 84.33495, 86.44958, 86.49708, 
    86.44078, 86.71569, 87.05787, 87.51586, 88.34952, 89.72784, 91.21667, 
    91.11954, 90.79993, 90.81182, 91.4836, 91.75092, 90.81039,
  86.42906, 85.2395, 84.68841, 84.98979, 84.85386, 83.55852, 81.75185, 
    81.728, 83.26623, 84.0872, 84.42953, 85.40857, 87.61354, 90.59848, 
    92.84652, 93.50609, 93.70979, 94.10858, 94.03317, 92.73042,
  90.10467, 88.99644, 87.46127, 84.8843, 80.96181, 77.44679, 75.36013, 
    74.95149, 76.64816, 78.92027, 81.20428, 83.4878, 86.1662, 89.42454, 
    92.43795, 93.59103, 92.74741, 92.09168, 92.38637, 92.77847,
  88.29583, 87.06824, 84.75077, 81.86219, 78.43339, 75.17641, 73.44144, 
    73.49783, 75.83514, 78.91843, 82.15327, 84.40033, 86.50436, 88.96901, 
    90.24062, 90.81704, 90.40244, 89.91724, 90.55677, 92.19358,
  85.10093, 82.53342, 78.77259, 75.51148, 73.2529, 72.13295, 72.46906, 
    74.07301, 77.45193, 80.78904, 83.28994, 84.61494, 85.96581, 87.69746, 
    88.53777, 88.77151, 88.70559, 88.65051, 89.92344, 90.82498,
  78.91714, 75.8001, 72.90591, 71.2389, 71.10546, 71.2846, 72.39175, 
    74.25391, 76.61257, 78.87014, 80.38984, 81.52134, 82.76875, 84.27552, 
    84.82957, 84.79922, 84.37336, 84.09708, 84.30559, 84.24113,
  74.92882, 72.61801, 71.87159, 72.0817, 72.55474, 72.29814, 71.73359, 
    69.43429, 66.27986, 66.35728, 68.52521, 72.21919, 75.80283, 77.49962, 
    78.69512, 79.52193, 78.63184, 76.78963, 76.29683, 77.17324,
  75.0826, 74.99387, 75.38715, 74.58057, 73.72732, 72.10017, 67.93317, 
    61.90069, 58.14434, 58.03096, 59.16175, 62.39209, 67.05926, 70.42199, 
    72.5098, 73.77815, 73.65945, 73.04981, 74.66146, 77.07867,
  72.18482, 71.63196, 69.91414, 68.15995, 67.40941, 66.29379, 64.02441, 
    59.88378, 58.57978, 60.45974, 60.71333, 62.75629, 67.49532, 71.65625, 
    74.12309, 74.77258, 74.58803, 74.62859, 75.61307, 76.20023,
  94.18742, 94.78651, 95.05796, 95.405, 95.78975, 96.09081, 95.82191, 
    96.29353, 95.64204, 95.16457, 95.92005, 96.58356, 96.23803, 96.38926, 
    97.45618, 97.08813, 96.43733, 97.22275, 97.09807, 96.88019,
  90.62778, 91.67963, 92.55199, 93.45461, 94.41479, 95.3639, 96.175, 
    96.91492, 93.30266, 93.83749, 94.09431, 94.44469, 95.0347, 95.58845, 
    95.99452, 97.05055, 95.33937, 96.01039, 96.49406, 97.16955,
  89.56061, 90.99419, 92.17153, 93.33259, 94.20679, 95.06, 95.84649, 
    96.58688, 92.36536, 93.25999, 94.1283, 94.91502, 95.64646, 96.33486, 
    96.89198, 97.33029, 96.19186, 97.22997, 97.79877, 98.45907,
  87.37453, 88.97194, 90.17204, 91.38701, 92.42426, 93.66591, 94.43172, 
    95.0938, 92.76897, 93.37857, 93.93302, 94.70012, 95.7581, 96.83466, 
    97.91909, 98.66738, 99.14138, 99.3316, 99.42347, 99.5379,
  84.02663, 85.7617, 87.41296, 88.39972, 88.76104, 89.11695, 89.75389, 
    90.31902, 89.81747, 90.62682, 91.36382, 92.09742, 92.75951, 93.36055, 
    93.78522, 94.57132, 97.65337, 97.66934, 97.57734, 97.56347,
  82.1002, 84.60815, 86.52597, 87.68933, 88.53323, 89.03803, 89.46874, 
    90.1379, 86.30141, 86.21947, 86.56834, 87.49635, 87.92371, 88.45892, 
    88.63931, 89.41075, 96.66512, 97.0029, 97.06432, 95.82013,
  88.79765, 87.70201, 88.24398, 88.81107, 89.85501, 91.0166, 90.36971, 
    89.45029, 80.87035, 79.59048, 78.43405, 75.60263, 76.20267, 81.00632, 
    84.68274, 80.13408, 87.65636, 91.09661, 93.63106, 94.56118,
  67.40107, 66.3269, 65.77606, 65.57142, 66.87114, 67.60163, 66.20417, 
    64.58878, 58.44157, 58.51526, 60.67277, 71.46075, 75.7475, 81.9043, 
    85.4471, 86.02991, 88.36167, 87.4909, 85.11867, 85.46948,
  80.07499, 78.7049, 78.11797, 78.20322, 78.35344, 78.12115, 77.83586, 
    76.94158, 74.4636, 73.96026, 73.65913, 74.07961, 76.4464, 79.39479, 
    79.95641, 79.73466, 80.26591, 82.15359, 84.80243, 87.83468,
  82.5872, 82.64403, 82.73331, 82.33069, 82.04414, 81.79884, 81.48571, 
    80.98991, 80.5477, 79.29243, 78.8994, 79.41393, 80.62057, 82.01878, 
    83.27122, 83.94476, 84.60968, 85.05183, 84.68274, 83.54757,
  82.30101, 82.36032, 82.1636, 82.30254, 82.55415, 82.4758, 82.0135, 
    81.55532, 81.53415, 80.97189, 80.97336, 82.02923, 83.29785, 84.32027, 
    84.53857, 84.36301, 85.07761, 86.4818, 87.84478, 87.70183,
  83.24864, 82.63571, 81.64894, 81.3427, 81.65742, 82.42092, 82.84842, 
    82.73674, 82.50926, 81.75832, 81.1097, 81.60217, 83.594, 85.88155, 
    86.80522, 86.55529, 86.92948, 87.88882, 89.15066, 89.00926,
  84.22817, 83.80845, 83.05275, 82.34894, 81.48191, 80.74599, 80.23893, 
    80.42862, 80.31598, 78.70084, 76.80389, 76.85663, 79.2311, 83.67585, 
    87.39967, 88.99288, 89.64552, 90.48902, 91.84641, 92.19759,
  85.04573, 84.55202, 83.81132, 81.83911, 78.25542, 75.35136, 73.67889, 
    73.22824, 73.15976, 73.12093, 73.35497, 74.95629, 77.98178, 82.19603, 
    86.12734, 88.16925, 88.96128, 90.11852, 91.59785, 92.2924,
  83.7087, 83.24825, 82.19896, 80.15905, 76.47398, 73.27189, 71.09848, 
    70.31129, 71.02663, 72.66221, 75.29576, 78.50362, 80.86558, 82.87668, 
    84.8227, 86.0659, 86.79785, 87.09083, 88.24793, 90.03617,
  81.48972, 80.61008, 78.42619, 75.52705, 72.63692, 71.03149, 70.82366, 
    71.84871, 73.92429, 76.71027, 79.49175, 81.48633, 82.36765, 83.24905, 
    84.11757, 84.50053, 84.44296, 84.35739, 85.98608, 87.6048,
  76.80487, 74.182, 72.01685, 70.96909, 70.85377, 71.33263, 72.83781, 
    74.49137, 75.95881, 77.74594, 79.16064, 80.25919, 80.98724, 81.79124, 
    82.25086, 82.15313, 82.01983, 81.77708, 82.18764, 83.23424,
  72.57234, 71.30907, 72.44624, 73.49619, 74.51273, 74.76886, 73.97821, 
    70.92802, 67.93851, 67.53635, 69.13773, 72.31934, 74.85915, 76.25638, 
    77.18455, 77.742, 77.5174, 76.79706, 77.07981, 77.73408,
  73.55667, 74.58836, 76.36998, 75.8345, 74.62085, 72.42974, 67.93636, 
    63.07016, 61.1617, 60.20385, 60.94213, 63.53188, 66.44196, 67.84573, 
    68.15906, 68.62862, 69.47968, 70.69564, 72.29819, 74.53253,
  72.17477, 72.20637, 71.11819, 70.63619, 70.4921, 68.50719, 66.60636, 
    63.37275, 62.90517, 62.44566, 60.69054, 62.0986, 65.4043, 67.15815, 
    67.07471, 67.4139, 68.68394, 70.88067, 73.07153, 74.40041,
  91.15734, 91.60645, 92.02863, 92.37306, 92.72182, 93.09782, 93.37084, 
    93.59296, 92.02976, 92.26305, 92.52608, 92.84922, 93.04916, 93.17595, 
    93.56516, 93.73692, 92.89298, 93.26173, 93.69658, 93.89421,
  84.89678, 86.26551, 87.77914, 89.36425, 90.93636, 92.48667, 93.85404, 
    94.96321, 91.84747, 92.54652, 92.8732, 93.24185, 93.69528, 94.17664, 
    94.87571, 95.39429, 94.06072, 94.836, 95.65474, 96.19641,
  83.33409, 85.633, 87.82729, 89.79224, 91.622, 93.11959, 94.08315, 94.9612, 
    91.09057, 92.49413, 93.22009, 94.08511, 94.79704, 94.29358, 94.63721, 
    94.87001, 93.9185, 94.82468, 95.90041, 96.95824,
  82.25124, 84.99084, 87.13528, 89.28705, 90.20464, 91.8223, 93.73186, 
    94.6946, 92.56321, 93.43413, 94.95737, 96.28828, 97.52716, 98.50653, 
    98.92906, 99.30764, 99.25262, 99.35851, 99.50764, 99.17085,
  80.148, 83.22833, 85.06017, 85.83403, 86.57191, 87.44714, 88.30205, 
    89.11346, 89.0246, 90.17924, 91.15912, 92.29076, 93.50791, 94.55234, 
    95.97889, 97.34693, 99.45856, 99.46698, 99.3004, 98.91789,
  80.64086, 83.13128, 85.10098, 86.19941, 87.00945, 87.25569, 87.35531, 
    87.39864, 82.44392, 81.82154, 82.25107, 83.26851, 84.60762, 86.06002, 
    87.08781, 87.61829, 93.98598, 94.8945, 95.81725, 96.01026,
  94.42855, 91.78777, 91.508, 91.22969, 90.49005, 90.45111, 89.89825, 
    90.2805, 83.02515, 83.81022, 84.56362, 75.24809, 76.08333, 80.64908, 
    85.64323, 80.4324, 86.9063, 89.59538, 91.93086, 93.4304,
  79.69307, 79.05977, 77.21204, 76.65639, 78.05148, 81.86672, 84.23633, 
    86.12074, 80.0108, 80.23608, 83.35241, 81.56915, 82.27223, 86.71738, 
    93.61224, 94.47672, 94.86639, 89.41753, 88.5628, 88.75526,
  68.86478, 66.18509, 63.97089, 62.28399, 61.3599, 61.14331, 60.70528, 
    60.10493, 57.95488, 58.09105, 60.57862, 66.33405, 71.72011, 76.58452, 
    78.72877, 80.92087, 85.2175, 90.46526, 94.12693, 94.52856,
  74.83242, 74.1268, 73.55509, 72.50199, 71.61811, 71.13254, 70.89545, 
    70.66103, 70.68108, 70.47277, 70.43621, 70.37753, 70.44761, 70.49295, 
    70.06162, 69.99065, 71.15992, 72.72083, 74.13442, 75.08565,
  79.46628, 79.07218, 78.22723, 77.53532, 77.39489, 76.79573, 76.01915, 
    75.16807, 74.67652, 74.35712, 74.38629, 75.14704, 76.05479, 76.88708, 
    77.50642, 77.88445, 78.4121, 79.10541, 80.10255, 80.78116,
  82.09145, 81.7422, 80.9482, 80.71723, 81.15379, 81.05611, 80.30183, 79.574, 
    78.58341, 77.39236, 76.28782, 76.36651, 77.7426, 79.31573, 80.27455, 
    80.61893, 80.97623, 81.81136, 82.88186, 83.48132,
  83.93591, 83.27991, 83.07052, 83.30554, 83.49915, 82.44849, 80.64565, 
    80.01933, 79.43593, 77.75064, 75.57474, 74.4676, 74.92387, 77.19232, 
    80.55775, 82.60503, 83.41345, 83.92077, 84.29457, 83.95155,
  86.93548, 86.24494, 85.89677, 84.94781, 82.5918, 79.93192, 77.60565, 
    76.35489, 75.60748, 75.21935, 74.56561, 74.6105, 76.21035, 79.25741, 
    82.45056, 84.32378, 84.23357, 84.03029, 84.22984, 84.58914,
  88.91182, 88.64409, 87.44064, 84.96096, 80.99002, 77.58259, 75.28165, 
    74.12822, 73.68913, 74.52712, 76.08347, 78.09045, 80.87344, 82.76668, 
    83.09406, 82.69834, 81.43202, 80.64182, 81.2855, 82.99592,
  85.88342, 85.78923, 83.31765, 79.49268, 75.78366, 73.82383, 73.37409, 
    73.88597, 74.99024, 77.31811, 80.23452, 82.99772, 84.31554, 83.70946, 
    81.48959, 79.78174, 77.84951, 76.74753, 77.74062, 79.14745,
  80.32345, 78.96923, 76.35722, 74.47417, 74.83141, 75.88432, 76.69282, 
    77.26063, 77.84904, 79.36651, 81.6597, 83.44891, 83.65135, 82.44675, 
    80.64413, 79.09695, 77.01386, 74.72459, 73.11312, 72.03884,
  78.15393, 76.33631, 76.97706, 78.70842, 80.61084, 81.17062, 79.06895, 
    73.00419, 67.21976, 65.53294, 67.66468, 70.984, 73.15779, 73.89642, 
    74.69585, 74.51506, 71.98235, 68.44883, 66.36206, 65.229,
  76.53444, 78.74321, 81.40226, 82.09846, 81.30482, 78.64753, 72.28579, 
    65.12807, 61.2155, 59.00515, 58.25527, 58.83998, 60.7355, 63.13327, 
    64.87085, 65.22993, 64.77605, 64.67072, 64.88647, 65.64855,
  72.93227, 74.04498, 74.42889, 74.49993, 74.65531, 73.2572, 70.20907, 
    65.31041, 64.99466, 65.15518, 61.02635, 59.48115, 62.1367, 64.85059, 
    65.27641, 65.55321, 66.02945, 66.99364, 68.12939, 68.67649,
  93.65504, 94.01929, 94.35616, 94.7345, 95.38509, 95.52082, 95.78677, 
    96.28745, 94.90966, 95.37086, 95.66442, 95.96046, 96.28737, 96.42122, 
    96.26952, 96.49857, 95.84058, 95.64158, 95.8696, 96.08067,
  88.48222, 89.74146, 90.95013, 92.43302, 93.81982, 95.21719, 96.30212, 
    97.1283, 93.96214, 94.70991, 95.23365, 95.70934, 96.23575, 96.85564, 
    97.68211, 98.2012, 97.04456, 97.62482, 97.55606, 98.20499,
  87.71947, 89.82251, 91.55999, 92.83865, 94.35081, 95.88737, 96.78246, 
    97.11669, 92.50648, 93.32105, 94.86143, 96.96326, 98.20955, 98.66987, 
    98.92329, 98.9958, 98.04813, 98.54354, 98.92281, 99.14491,
  88.50604, 90.20785, 91.40582, 92.46552, 93.43274, 94.14966, 95.54662, 
    96.49686, 95.36455, 96.8394, 97.57829, 97.77673, 97.98138, 98.79185, 
    99.39751, 99.60592, 99.90369, 99.94912, 99.9804, 99.98407,
  86.38065, 88.23083, 88.46715, 88.9861, 89.31184, 90.12469, 91.48721, 
    93.0732, 93.37662, 94.0401, 94.56462, 95.02261, 95.74331, 96.26222, 
    96.64214, 97.5881, 99.40902, 99.74716, 99.79674, 99.8482,
  86.57601, 88.11902, 89.33299, 89.50333, 90.27208, 90.48817, 91.4436, 
    92.55013, 88.64322, 89.18916, 89.80016, 90.47688, 91.25591, 92.30432, 
    93.35534, 94.39906, 98.87218, 99.13432, 99.22832, 98.80463,
  96.19411, 93.86968, 92.6435, 92.04849, 90.62171, 89.65601, 89.3793, 
    89.42174, 81.24668, 81.7877, 83.39718, 78.67282, 80.3922, 84.93423, 
    88.67194, 87.89617, 95.25839, 97.23863, 97.34412, 96.2718,
  95.71352, 94.65591, 92.80133, 91.34591, 91.99192, 92.9209, 93.69693, 
    93.86375, 86.6246, 86.98383, 88.35616, 84.22696, 84.06124, 89.05125, 
    92.25842, 94.34904, 96.19179, 96.6143, 93.72277, 94.127,
  80.42094, 80.44828, 81.78617, 82.80648, 83.48298, 83.41563, 82.87254, 
    81.44496, 79.71256, 81.95229, 86.51395, 89.48201, 90.89942, 91.71382, 
    90.89168, 90.29945, 92.10329, 94.41477, 95.35806, 95.18386,
  67.74119, 70.77429, 73.57495, 75.43352, 75.26719, 73.08345, 70.94035, 
    68.45725, 66.90898, 67.14294, 68.90697, 70.81448, 72.74093, 73.69423, 
    72.81675, 72.41267, 73.73449, 76.53379, 80.84863, 82.28402,
  69.0064, 69.59544, 69.23852, 69.20354, 68.68546, 66.92447, 66.18528, 
    66.58141, 68.25378, 70.16002, 72.70469, 75.39268, 77.40023, 78.83053, 
    79.34266, 79.24104, 79.09504, 78.29262, 76.98973, 74.4632,
  73.18201, 72.58765, 70.87976, 69.25682, 68.88557, 68.65481, 69.11671, 
    70.74843, 72.71302, 73.51521, 74.29568, 76.08853, 78.61827, 81.34708, 
    83.23657, 83.88277, 83.80129, 83.54655, 82.7213, 80.20423,
  75.28426, 74.78485, 73.66255, 72.69759, 72.72395, 71.93993, 70.70498, 
    70.88644, 72.0435, 72.34782, 72.42807, 72.89104, 74.36068, 77.21915, 
    81.14729, 84.08173, 84.52277, 84.1576, 83.58703, 82.43084,
  76.64052, 76.24683, 75.77996, 74.68929, 72.59476, 70.42841, 68.80214, 
    68.52505, 69.95641, 71.52836, 73.11008, 74.61452, 76.12936, 78.4775, 
    81.69926, 83.80149, 83.46873, 82.93182, 82.68647, 82.68516,
  77.28465, 76.68292, 75.40398, 72.82001, 68.68902, 65.5687, 64.33997, 
    65.67029, 68.89173, 72.129, 75.31797, 78.04042, 80.34892, 82.87875, 
    84.78902, 85.494, 84.56737, 82.92414, 81.90591, 81.79385,
  74.04151, 72.94321, 70.03185, 66.09653, 62.30177, 60.93573, 62.02865, 
    65.23481, 69.96077, 73.93886, 77.2197, 80.29555, 83.15405, 85.2132, 
    85.57269, 84.75986, 83.17626, 81.24062, 80.55569, 80.21854,
  70.27155, 67.4607, 63.92607, 61.26208, 60.77069, 62.78344, 65.83708, 
    69.09134, 72.49689, 75.13664, 78.00196, 80.81332, 83.04522, 84.14268, 
    83.9715, 83.34923, 81.62184, 79.06306, 76.77286, 75.16313,
  66.54787, 63.90538, 64.21473, 66.15341, 68.38175, 70.12006, 69.41013, 
    65.33405, 61.50743, 61.22532, 64.31711, 69.14079, 74.01866, 76.93654, 
    78.13708, 78.28484, 76.0531, 72.78801, 70.58049, 70.51802,
  65.69419, 66.74789, 68.99513, 69.72978, 69.3315, 66.10223, 60.5177, 
    55.71837, 54.02144, 53.01939, 53.53496, 55.92409, 60.67567, 66.21429, 
    69.76015, 71.2353, 71.18648, 70.87862, 71.09346, 72.42747,
  65.38427, 66.25015, 65.83321, 64.75883, 64.2741, 63.14878, 62.04262, 
    61.85006, 60.72356, 58.63106, 53.88764, 54.49686, 61.72274, 69.61214, 
    72.8765, 73.44109, 74.03866, 74.62927, 75.13474, 75.46233,
  90.80833, 91.20017, 91.56627, 92.12254, 92.60011, 93.05394, 93.45878, 
    93.83282, 92.67487, 93.21812, 93.59498, 93.89619, 94.31508, 94.60715, 
    94.92164, 95.29206, 94.72443, 95.06561, 95.15273, 95.02525,
  83.24882, 84.90469, 86.39455, 88.10995, 89.56744, 91.06527, 92.67813, 
    94.514, 91.55436, 92.74826, 93.63358, 94.24391, 94.89915, 95.6613, 
    96.50361, 97.26011, 95.92193, 97.00983, 97.62983, 98.14443,
  86.54725, 88.06969, 89.47744, 90.86056, 91.91708, 93.35291, 94.82675, 
    95.43842, 91.22856, 92.65474, 94.13358, 95.12713, 96.09125, 96.93686, 
    97.63849, 97.80606, 97.34197, 97.72067, 97.96343, 98.17055,
  86.48869, 88.00596, 90.0195, 91.60497, 92.95155, 94.35143, 95.70451, 
    96.99287, 96.55173, 97.23428, 97.29815, 97.69321, 98.08224, 98.33317, 
    98.50294, 98.48691, 98.63695, 98.66928, 98.7514, 98.90651,
  82.14108, 84.37273, 87.03036, 89.17256, 91.31558, 93.14911, 95.15055, 
    96.46055, 96.98433, 97.42814, 97.57892, 98.07599, 98.20596, 98.47234, 
    98.75258, 98.76122, 99.88519, 99.80664, 99.59342, 99.36972,
  80.60906, 82.4681, 85.02419, 87.52157, 89.44544, 90.96101, 92.05782, 
    92.61372, 88.38093, 88.93065, 89.82085, 91.00826, 92.30574, 93.73225, 
    95.13015, 95.98069, 99.533, 99.63696, 99.61808, 99.33809,
  92.59921, 89.15463, 88.47984, 89.09036, 89.48801, 89.92383, 89.93216, 
    89.76627, 81.78973, 82.87427, 85.28613, 82.25102, 84.35693, 91.20017, 
    92.03934, 91.30197, 95.33393, 95.96706, 96.1652, 95.96898,
  95.69055, 95.32285, 95.32874, 95.83955, 96.29237, 96.87567, 97.29719, 
    97.77764, 95.68285, 96.05286, 96.79561, 94.7751, 93.89149, 95.35786, 
    95.51825, 96.31172, 96.94995, 97.17868, 95.13857, 95.43344,
  97.56347, 97.09823, 95.66154, 95.69984, 96.82388, 97.89753, 98.77161, 
    98.88055, 97.0269, 97.09394, 97.47529, 97.48767, 97.19893, 96.93158, 
    96.44757, 96.54613, 97.47803, 98.04446, 97.98174, 97.25314,
  97.6192, 97.29438, 96.81134, 96.53033, 96.8, 96.2001, 96.21688, 96.67461, 
    96.99799, 96.05125, 93.94894, 92.57611, 92.1538, 91.90034, 91.44589, 
    90.13371, 91.13171, 93.40109, 95.15395, 95.11039,
  84.84947, 85.2535, 86.62653, 89.43372, 90.91171, 89.62801, 88.47688, 
    87.38583, 85.48166, 80.5733, 76.21326, 74.72947, 74.04553, 73.18244, 
    72.97602, 71.39422, 70.66349, 71.45934, 73.86978, 74.91567,
  67.46163, 68.24608, 69.17294, 70.2288, 70.37189, 69.42071, 68.23119, 
    67.85434, 67.67406, 66.27837, 65.08662, 64.95678, 66.32552, 68.63753, 
    70.76314, 72.00292, 72.48904, 73.17322, 73.89768, 73.99493,
  68.96284, 69.54314, 69.86569, 69.77566, 68.90533, 67.04539, 64.98909, 
    64.32863, 64.87811, 65.17906, 64.95242, 65.07683, 66.17075, 68.69654, 
    73.24338, 76.85174, 78.36485, 79.21473, 79.54841, 78.85603,
  71.68563, 71.50587, 71.47861, 70.95265, 69.39536, 67.3045, 65.47205, 
    64.99845, 66.24803, 68.30613, 69.91898, 71.59579, 72.85583, 74.42352, 
    77.35901, 79.47066, 79.99783, 80.293, 80.57137, 80.65427,
  72.12289, 72.51076, 72.61028, 71.67716, 68.69285, 66.01337, 63.89356, 
    63.913, 66.44003, 70.4908, 73.87232, 76.31756, 77.83153, 78.9334, 
    80.26783, 81.10192, 80.80811, 79.86362, 79.83588, 80.94078,
  72.8618, 73.2907, 71.97399, 68.63506, 64.72836, 62.98349, 63.26275, 
    65.71283, 70.25196, 74.70642, 77.70745, 79.75386, 80.98125, 82.22801, 
    82.85043, 82.24965, 80.47363, 78.50451, 78.65433, 79.50929,
  69.7233, 67.98829, 64.87098, 62.15294, 61.63873, 63.67168, 67.34159, 
    71.38271, 74.8109, 76.99274, 78.87776, 80.57784, 81.83745, 82.83095, 
    82.42424, 81.26121, 79.10313, 76.73915, 75.03993, 73.98985,
  65.71285, 63.70486, 64.07835, 66.67607, 69.88301, 73.19782, 74.0668, 
    70.89298, 66.86757, 65.70147, 67.13364, 70.46742, 74.1769, 76.08712, 
    77.30626, 77.70287, 74.61949, 70.9513, 69.07899, 68.45926,
  68.75172, 71.02628, 74.31329, 76.97478, 77.42233, 73.70608, 67.11523, 
    61.20573, 57.99365, 55.24018, 53.99352, 55.36421, 59.22341, 63.63469, 
    66.68666, 68.15988, 67.78951, 66.9177, 67.08877, 67.50816,
  71.92353, 74.6707, 76.11405, 76.31284, 74.72383, 70.79923, 67.66563, 
    66.98893, 65.3332, 63.40308, 56.91211, 55.98566, 61.25433, 67.31401, 
    69.73647, 70.42716, 70.84703, 71.37173, 71.90376, 71.7758,
  93.19692, 93.10423, 93.5722, 94.34063, 94.46259, 94.81142, 95.19144, 
    95.45174, 94.20775, 94.84272, 95.1311, 95.02566, 95.84089, 96.15184, 
    96.46856, 96.80448, 96.02759, 96.69588, 96.69997, 96.87078,
  86.93295, 88.29019, 89.70782, 90.87581, 92.17657, 93.27828, 94.28043, 
    95.50006, 92.19778, 92.70957, 93.41745, 94.59193, 95.33624, 96.11549, 
    96.37658, 96.91048, 95.22714, 96.34199, 96.51436, 97.36287,
  85.47877, 87.1825, 89.21128, 91.31468, 93.03142, 94.17542, 94.90562, 
    95.80197, 91.06454, 92.27455, 93.41293, 94.61885, 96.01, 97.12698, 
    98.17449, 98.64558, 98.06181, 98.58057, 98.5295, 98.55048,
  84.81056, 86.72003, 89.23831, 91.54677, 93.26199, 94.35738, 95.41176, 
    96.44925, 95.07298, 97.09825, 98.55858, 99.15589, 99.65255, 99.77599, 
    99.8498, 99.82594, 99.75752, 99.59941, 99.38647, 99.1387,
  83.43355, 86.52654, 88.80086, 90.39192, 91.15159, 92.40733, 94.05563, 
    95.6782, 96.29297, 97.546, 97.57794, 96.71319, 96.79937, 96.80756, 
    96.86359, 97.28355, 99.06136, 99.30521, 99.1705, 99.18734,
  80.44089, 83.43877, 85.30309, 86.00222, 86.06197, 86.76756, 87.76027, 
    88.78304, 85.19894, 85.42948, 85.72399, 85.64291, 86.6544, 87.40753, 
    88.53481, 90.03323, 96.59608, 97.61682, 98.07783, 97.8933,
  97.16106, 92.73128, 92.69839, 91.1569, 89.70806, 88.93984, 88.80118, 
    88.6536, 80.73916, 81.01459, 83.15285, 75.85268, 77.82914, 85.37975, 
    86.32574, 81.85006, 88.77656, 91.35705, 92.90398, 93.5135,
  99.50124, 99.28654, 97.91061, 96.10656, 95.34344, 95.48924, 95.48679, 
    95.47013, 92.32063, 94.10294, 96.99541, 93.43474, 94.30569, 97.42249, 
    97.14465, 94.91272, 95.49815, 95.28429, 86.22903, 85.84734,
  97.90517, 98.23191, 98.39751, 98.12723, 98.40765, 98.44724, 98.16487, 
    97.98857, 95.80811, 96.02682, 97.13729, 97.79931, 97.80248, 97.40653, 
    97.27087, 97.99877, 98.3995, 99.27049, 99.11123, 98.98117,
  97.47858, 97.09048, 96.65763, 96.68069, 96.57857, 96.26048, 96.19877, 
    96.18422, 96.23477, 96.17944, 96.34633, 96.98767, 97.81219, 98.21944, 
    98.63589, 99.06728, 99.05439, 98.92059, 98.53691, 97.80628,
  96.57491, 96.12096, 96.13557, 95.82262, 95.96558, 95.64795, 95.3382, 
    94.81771, 93.81004, 92.0926, 90.6209, 89.59002, 90.07716, 91.82098, 
    93.25934, 93.65376, 93.78416, 94.09309, 94.10136, 95.03428,
  87.74431, 87.14758, 86.70133, 86.74864, 87.17286, 84.69859, 78.95452, 
    75.66056, 71.61276, 66.62209, 63.38577, 62.07311, 63.24553, 66.7522, 
    69.98003, 71.50812, 73.43144, 76.71527, 78.67895, 74.00208,
  71.97076, 70.67438, 69.61774, 69.28181, 68.9511, 68.0744, 66.34554, 
    66.04761, 66.57143, 65.92511, 64.65747, 64.17191, 64.54499, 66.46928, 
    69.98008, 72.77322, 73.43833, 73.14802, 72.1029, 69.722,
  72.72495, 73.16222, 73.41911, 72.3142, 69.7308, 67.47719, 66.09325, 
    65.97969, 67.27386, 69.19496, 70.5024, 71.38602, 72.59468, 74.18335, 
    76.80907, 79.1534, 79.32914, 79.25886, 79.36954, 78.98549,
  74.74873, 75.15179, 74.87167, 73.34528, 69.60639, 66.57464, 64.41036, 
    63.97453, 66.1374, 69.75564, 73.32148, 76.25613, 78.47682, 79.61513, 
    80.6607, 81.77293, 81.88025, 81.13052, 81.07678, 82.08966,
  73.41413, 73.01344, 70.88447, 67.36964, 63.38716, 61.44658, 61.42782, 
    63.55565, 68.22065, 73.97116, 78.73363, 81.76145, 83.59144, 85.08396, 
    86.01371, 86.08192, 84.83362, 82.63183, 81.89792, 82.14648,
  69.18513, 65.61463, 60.97953, 57.58144, 56.28502, 57.5615, 60.43177, 
    64.69913, 70.07455, 74.80454, 78.55631, 81.82968, 84.04293, 85.49791, 
    86.22974, 86.09874, 84.41599, 81.99628, 79.61255, 77.77396,
  62.1845, 57.94397, 56.86998, 58.0495, 60.79956, 64.69273, 67.83666, 
    67.04001, 64.51396, 63.85782, 66.74741, 71.96326, 76.27963, 78.50108, 
    79.99211, 80.51544, 78.48409, 74.85291, 71.82368, 70.36896,
  63.10419, 63.74438, 65.86459, 68.9133, 71.07522, 69.30617, 64.37768, 
    59.822, 57.93431, 55.55207, 55.71085, 58.76806, 63.2041, 66.105, 
    67.15285, 67.35664, 66.34543, 65.26459, 65.05976, 65.66129,
  67.66135, 68.30825, 68.40594, 68.66152, 66.797, 63.27365, 61.69573, 
    63.57627, 64.04705, 62.19039, 57.6351, 57.87633, 63.19652, 66.07482, 
    65.58461, 65.44444, 66.1988, 67.17632, 67.67261, 68.33199,
  89.97185, 90.5379, 90.8612, 91.38109, 91.72076, 92.19814, 92.60293, 
    92.98607, 91.91235, 92.41994, 92.87119, 93.3403, 93.77194, 94.05481, 
    94.31158, 94.452, 93.75748, 93.8994, 93.95657, 93.89941,
  83.7226, 85.47976, 87.28371, 89.13623, 90.7288, 92.10673, 93.18844, 
    93.99819, 90.35492, 91.51194, 92.35429, 93.07935, 93.76382, 94.53299, 
    95.86916, 96.4803, 95.13585, 96.33618, 97.33565, 97.95048,
  86.84631, 89.02713, 90.91268, 92.46983, 93.92436, 95.03396, 95.38171, 
    95.57854, 91.14893, 92.61815, 93.89426, 95.47335, 96.90436, 97.85351, 
    98.38326, 98.76429, 98.18401, 98.69257, 98.89284, 99.20484,
  87.87009, 89.55447, 90.33923, 91.43469, 92.67441, 94.21761, 95.51057, 
    96.18581, 94.30418, 94.71414, 95.03587, 95.49099, 97.00898, 98.27115, 
    99.14165, 99.39479, 99.10202, 98.94683, 98.41821, 97.59863,
  86.04722, 88.76143, 89.99367, 90.34675, 90.91614, 91.16277, 91.54984, 
    92.00558, 90.34175, 90.66476, 92.30382, 93.70452, 95.09856, 96.6235, 
    97.59767, 97.85804, 99.05326, 98.97215, 98.20609, 97.87965,
  82.81487, 84.13323, 84.54802, 84.15417, 83.96962, 83.97035, 83.42916, 
    84.12977, 80.11827, 81.54885, 83.64851, 85.50327, 86.96062, 88.40745, 
    89.80241, 91.85929, 97.23978, 97.97952, 98.5767, 98.34953,
  93.40611, 90.46309, 89.73368, 88.3972, 86.48867, 85.23512, 83.70213, 
    82.14357, 74.10271, 75.00026, 78.12263, 70.04846, 71.54284, 80.84724, 
    83.06602, 79.72066, 88.84737, 91.68056, 93.41286, 94.51488,
  96.35163, 95.99653, 95.42265, 94.55402, 94.16482, 94.03839, 94.38236, 
    95.03768, 91.63159, 92.31866, 93.83195, 92.5961, 92.07475, 94.97099, 
    95.87269, 88.76534, 92.97592, 92.02648, 88.37914, 90.77307,
  98.19268, 98.46968, 98.42301, 98.08195, 97.75488, 97.2318, 96.28963, 
    95.19823, 93.137, 94.1226, 95.77103, 96.72723, 96.6893, 95.97787, 
    95.53902, 95.82535, 96.76891, 98.08115, 98.10097, 98.04954,
  97.18988, 97.24141, 97.28095, 97.58509, 97.50785, 97.34171, 96.70387, 
    96.05, 95.13084, 94.68771, 95.08193, 95.9284, 96.32025, 95.81417, 
    95.81268, 95.90349, 95.77541, 96.60865, 97.21698, 97.18893,
  96.18966, 96.28281, 96.13585, 96.02641, 95.71938, 95.85464, 95.937, 
    96.06284, 96.06138, 96.17554, 96.18291, 95.5539, 94.13596, 92.96144, 
    93.59525, 94.62584, 94.53702, 94.45964, 94.14228, 94.70921,
  93.56349, 93.53648, 93.63116, 92.85789, 93.2752, 93.0766, 92.9112, 
    92.68549, 91.01975, 87.46516, 82.8755, 76.24386, 72.82621, 74.67329, 
    80.82408, 89.03349, 90.65365, 91.14637, 91.09148, 91.47551,
  86.2842, 84.27705, 83.19467, 80.89996, 79.93822, 77.07063, 73.92938, 
    72.79076, 71.67305, 69.27796, 66.51881, 64.90306, 64.1787, 64.18735, 
    65.38896, 67.09972, 68.23392, 69.693, 70.8717, 69.54637,
  79.97189, 79.22208, 78.49727, 77.23862, 75.26921, 73.14004, 71.65726, 
    71.09402, 70.79529, 70.58079, 69.60879, 69.01481, 69.18788, 69.79019, 
    70.3418, 71.03977, 70.25855, 69.88831, 69.98515, 69.92155,
  81.01139, 81.03554, 79.88729, 77.70427, 74.43412, 71.80734, 69.79896, 
    68.75513, 69.27589, 70.52196, 71.55629, 72.70222, 73.9284, 74.53105, 
    74.45898, 74.46779, 73.76376, 72.87569, 73.04027, 74.55908,
  82.16694, 81.66604, 78.96965, 75.02692, 71.18566, 69.20417, 68.40496, 
    68.82653, 70.81581, 73.72656, 76.24717, 77.79568, 78.55941, 78.76706, 
    78.4638, 78.03761, 76.4044, 74.42401, 73.83415, 74.47393,
  82.21838, 79.37792, 75.06048, 70.92255, 68.76475, 68.71758, 69.68054, 
    71.09093, 73.39808, 75.30704, 76.75883, 78.07467, 79.08884, 79.91271, 
    79.59512, 78.54958, 76.15627, 73.52505, 71.04167, 69.0561,
  77.54633, 72.57208, 70.89728, 71.1451, 72.37165, 74.20956, 75.23063, 
    71.51285, 66.62112, 65.05525, 66.23386, 68.65853, 71.03112, 72.80261, 
    73.74546, 73.48061, 70.31933, 66.39304, 63.42192, 62.09817,
  74.18047, 74.89134, 75.85868, 75.75273, 75.91942, 74.40553, 69.59779, 
    63.91706, 60.75214, 57.44518, 56.61284, 57.71228, 60.18162, 61.83186, 
    63.32606, 64.52855, 64.44444, 63.96606, 63.55253, 63.60842,
  74.83121, 74.83449, 74.0708, 72.31294, 71.08938, 68.45897, 66.71553, 
    67.45971, 67.73402, 64.68311, 59.16714, 58.56633, 64.66608, 68.49735, 
    68.74585, 69.22419, 70.26541, 71.12468, 71.04853, 70.32848,
  93.35609, 93.79854, 94.24268, 94.59473, 95.0124, 95.22878, 95.49422, 
    95.83595, 94.56722, 94.85726, 95.02065, 95.27592, 95.90985, 96.49706, 
    96.79742, 96.82733, 96.13255, 96.2345, 96.85018, 97.13223,
  86.80276, 87.94537, 89.27338, 90.64491, 92.09734, 93.51076, 94.55887, 
    95.51414, 91.80738, 92.1687, 92.5789, 93.29871, 94.17729, 94.71819, 
    95.32184, 96.22286, 94.94872, 96.53972, 96.94118, 98.02116,
  85.43485, 87.50179, 89.40009, 91.02656, 92.33701, 93.57665, 94.6035, 
    95.57886, 91.66554, 92.85368, 93.34785, 94.46449, 95.6429, 96.57581, 
    97.40749, 97.86311, 97.51188, 97.9281, 98.12807, 98.54559,
  86.28155, 88.18664, 90.26792, 92.62183, 94.07873, 95.01184, 95.72089, 
    96.27785, 94.35239, 95.45249, 96.43911, 97.41747, 98.37515, 98.94194, 
    99.21447, 99.34201, 99.43716, 99.19517, 98.66732, 98.36206,
  82.8195, 84.4305, 86.4137, 87.60162, 88.43552, 89.70311, 90.68896, 
    91.74966, 92.00491, 93.17906, 94.22277, 94.93931, 95.30679, 95.76054, 
    96.21206, 96.27317, 98.34898, 98.51225, 98.92977, 98.90226,
  80.05388, 81.33138, 83.33538, 84.71581, 86.01432, 86.75815, 87.30588, 
    87.44364, 82.28201, 82.76255, 83.377, 83.73605, 84.92885, 85.90309, 
    86.70953, 87.75502, 94.46098, 96.02417, 96.9755, 96.61068,
  93.25208, 90.64008, 90.86642, 90.60185, 89.94553, 90.02608, 89.98444, 
    89.79893, 81.9163, 82.53802, 84.58971, 76.88049, 77.99996, 84.10915, 
    86.42484, 83.22768, 89.45352, 91.14999, 92.3505, 92.58658,
  97.16766, 97.21783, 97.42146, 97.43887, 98.13538, 98.17981, 98.30367, 
    98.49921, 93.51938, 94.33084, 94.90618, 91.58392, 91.74155, 95.40824, 
    97.19741, 87.53819, 94.76686, 92.32295, 88.52798, 88.66811,
  97.34184, 97.44157, 97.22591, 96.82339, 96.89909, 97.02335, 96.4408, 
    96.50729, 95.41898, 95.84706, 96.26937, 96.45774, 96.48514, 96.43723, 
    96.71026, 97.54182, 97.52422, 98.45792, 98.13587, 98.26196,
  96.08366, 95.89207, 95.80476, 95.90109, 96.05621, 95.94827, 96.03421, 
    95.96251, 95.86641, 96.31217, 96.86523, 97.29394, 97.35397, 97.14762, 
    96.78527, 96.96413, 97.10602, 97.14011, 96.8367, 96.43974,
  94.34266, 93.81937, 93.46854, 93.85558, 94.4488, 94.61611, 94.51689, 
    94.35003, 94.61697, 94.75643, 94.48959, 94.71329, 94.80341, 94.76806, 
    94.45033, 94.09579, 93.68062, 93.65158, 93.83111, 94.2262,
  93.98348, 93.63507, 93.21581, 92.75313, 92.54426, 92.55757, 92.25179, 
    91.98569, 91.31821, 88.80456, 84.60566, 81.51987, 80.26688, 81.28648, 
    86.82955, 89.03196, 88.79266, 88.37222, 88.87456, 89.41383,
  92.85101, 92.37439, 91.40523, 90.06389, 86.51424, 83.17644, 77.79111, 
    74.35162, 73.48146, 71.92123, 69.40263, 68.02954, 68.43786, 70.10921, 
    72.64298, 75.20477, 76.37994, 77.10701, 77.73832, 77.38582,
  81.4097, 80.53878, 79.04382, 77.24047, 74.51345, 71.96215, 70.04441, 
    69.63322, 70.71638, 72.07213, 72.39566, 72.77956, 74.13577, 75.92496, 
    77.1255, 77.89571, 77.68119, 77.5254, 77.66862, 77.66991,
  80.78194, 80.85741, 79.89391, 77.74844, 74.10768, 71.29113, 69.4744, 
    69.15372, 70.66894, 72.83791, 75.08286, 77.4659, 79.48566, 80.84589, 
    80.73795, 80.39294, 80.08677, 79.77051, 80.07536, 81.95976,
  79.55669, 79.52367, 77.31916, 72.97009, 68.15695, 66.0257, 65.79095, 
    66.86116, 69.69061, 73.55396, 77.80607, 80.74821, 82.5611, 83.32446, 
    83.0182, 83.09333, 83.00255, 82.03437, 81.94509, 83.35925,
  75.84201, 73.01212, 68.7271, 64.76467, 62.37858, 62.84763, 64.56116, 
    66.75629, 70.05988, 73.94013, 77.42159, 80.11255, 81.95464, 82.87777, 
    82.46145, 82.30193, 81.20995, 79.65732, 78.17568, 77.19614,
  68.80405, 64.45102, 62.9844, 63.27937, 64.56976, 67.09783, 69.56747, 
    68.12286, 65.09658, 64.95383, 66.92312, 70.12794, 73.71107, 75.61591, 
    76.64703, 76.70284, 74.31042, 70.89841, 68.0921, 66.26343,
  66.53922, 66.99717, 68.48034, 70.27734, 72.14618, 71.49644, 66.89308, 
    62.06602, 60.00855, 57.21362, 55.34502, 56.62545, 59.59315, 61.82316, 
    63.23282, 63.55645, 62.16237, 60.66155, 60.21361, 60.67094,
  69.7756, 70.76102, 71.48158, 70.62247, 68.29648, 65.12076, 63.44077, 
    63.60076, 63.64088, 60.32219, 56.42892, 56.07934, 61.38632, 64.29739, 
    64.70737, 64.39137, 63.47762, 63.09828, 63.6133, 65.21372,
  87.87144, 88.21857, 88.60684, 88.94148, 89.31792, 89.68599, 90.07487, 
    90.45275, 89.00296, 89.30055, 89.56355, 89.80946, 90.02379, 90.26151, 
    90.5332, 90.7392, 89.87868, 90.07836, 90.29291, 90.49884,
  80.42849, 81.60761, 82.88245, 84.32142, 85.68339, 87.12811, 88.41635, 
    89.99606, 87.29495, 88.6852, 90.019, 91.64638, 93.04214, 94.34138, 
    95.22759, 95.99899, 95.05128, 95.849, 96.43544, 96.83157,
  81.6123, 83.45866, 85.34392, 87.29916, 88.99227, 90.46492, 91.74153, 
    92.8705, 88.51039, 89.38605, 90.31899, 91.6171, 93.15782, 94.40815, 
    95.69617, 96.89381, 96.08431, 96.8004, 97.51286, 97.91598,
  85.27851, 86.83308, 88.48684, 90.12324, 91.41131, 92.47855, 93.78951, 
    95.19258, 92.98, 93.73174, 94.48363, 95.41576, 96.20052, 97.04327, 
    97.62795, 97.82314, 98.37493, 98.35964, 98.25789, 98.01603,
  83.99516, 86.16203, 88.64035, 90.977, 92.15356, 92.78673, 93.27843, 
    93.57978, 92.60374, 93.59895, 94.21228, 95.14954, 95.97317, 96.62777, 
    96.99928, 97.0396, 99.21751, 99.11832, 98.99919, 98.71571,
  83.11343, 84.92762, 86.26138, 87.49755, 87.91591, 87.46304, 87.12009, 
    87.30718, 83.25497, 83.58852, 84.27411, 85.43165, 86.70168, 87.78777, 
    89.06363, 90.40202, 97.01114, 97.56322, 97.51183, 96.42073,
  92.49075, 91.65252, 90.70885, 89.81654, 89.75542, 90.09502, 89.50841, 
    88.91155, 81.04165, 81.47257, 81.82097, 76.12496, 77.02622, 82.86564, 
    83.98397, 81.49069, 88.64997, 91.1809, 92.94584, 93.71318,
  95.32759, 95.4461, 94.77758, 93.9317, 94.24052, 94.72199, 95.36882, 
    95.62968, 91.49686, 91.46371, 89.7354, 87.81973, 89.34557, 93.18307, 
    94.68163, 85.35271, 92.37055, 90.4427, 86.9918, 88.62218,
  96.3307, 96.08435, 95.95122, 95.16783, 94.90248, 94.97745, 95.07863, 
    94.47644, 92.33926, 92.65597, 93.09394, 93.51646, 93.4259, 92.96649, 
    93.51923, 94.18346, 93.9185, 94.95898, 95.45123, 95.54339,
  95.2508, 95.29099, 95.34182, 95.68542, 96.11112, 95.96671, 95.61362, 
    95.04787, 95.08445, 94.95713, 95.00121, 95.42138, 95.2666, 94.69317, 
    94.75959, 94.52868, 94.04987, 93.84427, 94.27265, 93.94214,
  94.52175, 94.40124, 94.43031, 94.80775, 95.33078, 95.49467, 95.24235, 
    94.9965, 94.92789, 94.54887, 94.64713, 94.67353, 94.38345, 94.02478, 
    93.97343, 93.59296, 92.71645, 92.15865, 91.74821, 91.59586,
  95.2411, 94.77441, 94.04901, 93.4119, 93.54272, 94.11973, 94.16108, 
    93.67728, 92.86369, 91.69766, 89.46271, 87.4464, 87.09272, 87.27465, 
    89.05686, 90.21342, 90.38181, 90.29891, 90.59447, 90.67177,
  94.0123, 92.77683, 91.53129, 90.36688, 89.2187, 88.33691, 85.33851, 
    82.05627, 80.20957, 77.4863, 72.65121, 69.49371, 69.70012, 71.69787, 
    74.47786, 77.02297, 78.20784, 78.97698, 79.82038, 79.84093,
  87.65218, 85.5228, 83.29674, 80.86729, 78.14963, 75.6125, 73.48176, 
    72.26075, 71.68211, 72.03935, 71.81115, 71.93524, 73.07524, 75.07526, 
    76.76811, 77.54896, 77.39342, 77.86041, 78.99825, 80.21004,
  87.36882, 86.25879, 84.73042, 82.25171, 78.64264, 75.52785, 72.72984, 
    70.9302, 70.62196, 71.80356, 73.03072, 74.66441, 76.64874, 78.44851, 
    79.09248, 78.9557, 78.49244, 78.87772, 80.1887, 82.82592,
  87.26636, 86.56229, 84.17401, 79.85969, 74.9259, 72.3065, 71.11485, 
    70.9416, 71.6984, 73.62904, 76.12592, 78.66496, 80.68913, 81.76509, 
    81.12311, 80.60557, 80.21279, 79.6226, 79.70898, 81.11452,
  83.12348, 80.6437, 76.11108, 70.72128, 67.75606, 67.81651, 69.40057, 
    70.98038, 72.22362, 73.44923, 75.52654, 77.99159, 80.00219, 80.9564, 
    80.18394, 79.31335, 78.06211, 76.66676, 75.47005, 75.01969,
  74.94019, 69.92715, 67.75098, 67.01234, 67.70231, 69.55949, 71.20536, 
    68.85271, 64.65533, 63.45084, 64.95639, 68.12385, 71.65762, 73.83953, 
    74.75122, 74.50492, 72.60168, 70.21142, 68.69592, 67.71815,
  70.36284, 72.02059, 73.46619, 73.65868, 74.49564, 74.20656, 69.45376, 
    63.34934, 60.09494, 58.24009, 58.20577, 59.49382, 61.80649, 63.83165, 
    65.74013, 66.57152, 66.75034, 66.58237, 66.66656, 66.92596,
  72.15268, 73.95309, 74.01937, 74.45081, 74.13342, 72.31393, 68.99811, 
    65.39091, 64.90012, 62.41132, 60.1097, 61.04702, 66.21744, 68.95999, 
    69.49941, 69.88156, 70.08851, 70.16541, 70.60847, 71.22608,
  90.12871, 90.50231, 90.94535, 91.3054, 91.66551, 92.05522, 92.42523, 
    92.72335, 91.35476, 91.68061, 92.03687, 92.41409, 92.79233, 93.16836, 
    93.52808, 93.84317, 92.94817, 93.2752, 93.54611, 93.76267,
  84.33915, 85.03479, 85.93497, 86.86361, 87.72723, 88.61031, 89.672, 90.755, 
    87.54777, 88.34738, 89.23812, 90.26182, 91.41325, 92.35338, 93.37205, 
    94.18561, 92.49188, 93.4042, 94.13689, 94.72624,
  81.27549, 82.59588, 83.956, 85.57547, 87.24921, 88.75264, 90.04071, 
    91.24249, 86.92419, 87.90252, 88.7399, 89.75381, 90.91251, 91.96198, 
    93.30394, 94.76257, 93.61117, 94.47108, 95.06218, 95.66415,
  82.36783, 84.15694, 85.95633, 87.86015, 89.39191, 91.03252, 92.52575, 
    93.81688, 91.36697, 92.10178, 92.96253, 93.66862, 94.2865, 94.68461, 
    94.94682, 95.2058, 96.20732, 96.33025, 96.20891, 95.98954,
  82.44287, 84.94718, 87.1204, 88.66627, 90.21811, 91.06269, 92.05679, 
    93.08578, 92.31574, 92.9489, 93.23389, 93.79758, 94.29402, 94.60776, 
    94.77901, 95.06092, 98.7331, 98.48241, 98.02011, 97.53481,
  83.4572, 84.99305, 86.25269, 87.34988, 88.08547, 88.85759, 89.31202, 
    89.73009, 85.75915, 86.12881, 86.59358, 87.45907, 88.6804, 90.27583, 
    91.73309, 93.04957, 98.62062, 98.8606, 98.79662, 98.41615,
  90.86416, 88.93733, 87.3681, 87.33153, 87.26092, 87.62371, 87.81396, 88.14, 
    80.98979, 81.7655, 81.08409, 79.77519, 81.21045, 86.46884, 88.19651, 
    88.12832, 95.11156, 96.96672, 98.05554, 98.58126,
  94.46326, 94.42244, 94.02035, 94.06783, 93.78584, 93.80173, 94.18226, 
    94.23003, 89.98696, 89.88605, 85.47248, 86.53645, 87.83334, 91.96561, 
    92.04295, 80.89352, 89.32606, 95.33126, 95.86481, 97.31301,
  97.0152, 96.52802, 95.93153, 95.75603, 95.62247, 94.78349, 93.42371, 
    92.49545, 90.50257, 90.56016, 90.02274, 89.55293, 90.17064, 91.08939, 
    92.57377, 93.51434, 92.72825, 92.19247, 91.91468, 94.40428,
  96.52115, 96.68314, 96.65623, 96.30122, 96.45524, 96.43048, 96.20654, 
    95.97614, 95.52072, 95.29065, 94.61665, 94.15576, 93.6734, 93.29665, 
    93.64252, 94.26466, 94.4026, 94.55314, 94.92516, 95.32675,
  95.92165, 95.96313, 95.85695, 95.59916, 95.65395, 95.76101, 95.65024, 
    95.371, 94.94408, 94.62546, 94.2742, 94.2421, 94.43598, 94.24173, 
    93.70036, 93.60335, 93.08978, 92.89485, 93.07232, 93.19593,
  95.72863, 95.42015, 94.90595, 94.51858, 94.50774, 94.33872, 94.24818, 
    94.20869, 92.9856, 92.27758, 91.60546, 91.3122, 91.90127, 92.57652, 
    92.90247, 92.71616, 91.92661, 91.23918, 91.06407, 91.03968,
  91.45636, 91.0639, 90.75691, 90.29784, 89.31352, 87.76302, 85.25755, 
    84.36756, 83.52965, 81.65321, 77.88171, 75.33541, 76.30077, 79.01105, 
    80.64036, 81.8775, 82.23154, 82.7098, 83.66405, 84.68908,
  87.88451, 87.38002, 86.96318, 85.99594, 83.44963, 79.99928, 77.00716, 
    75.4815, 74.47584, 74.85666, 74.43276, 74.21986, 75.45686, 77.49866, 
    79.3102, 80.39404, 80.2767, 81.03935, 82.62309, 84.65954,
  86.6539, 86.60459, 85.85606, 83.54576, 79.52264, 75.76987, 72.36401, 
    70.12865, 69.42846, 70.76504, 72.42073, 74.26367, 76.4174, 78.1579, 
    79.19598, 79.72649, 79.50046, 80.20208, 82.22504, 85.29313,
  84.99163, 84.85098, 82.44604, 78.30439, 73.88101, 70.96342, 69.08198, 
    68.03592, 67.82262, 69.55432, 72.06441, 74.58332, 76.6958, 78.46339, 
    78.23687, 77.76344, 77.67222, 77.82519, 78.88546, 80.84192,
  82.77914, 81.13661, 77.3871, 73.12724, 70.7853, 70.09842, 69.63857, 
    68.9789, 68.39246, 69.11364, 70.53811, 72.52351, 74.44175, 75.92553, 
    75.52361, 74.23152, 72.43055, 70.91119, 70.02615, 70.15419,
  81.3384, 78.08202, 75.01406, 73.08229, 72.78662, 72.31483, 71.09338, 
    66.97353, 61.30368, 59.12077, 59.88459, 61.98553, 64.48939, 66.4251, 
    67.34624, 67.22649, 64.66857, 61.72177, 60.26021, 60.81456,
  79.63127, 78.33132, 77.04567, 76.09246, 75.69939, 73.14751, 67.77194, 
    62.00335, 56.09146, 52.82872, 51.96465, 53.33188, 55.68167, 57.46814, 
    58.6763, 59.24568, 58.76416, 58.4878, 59.51992, 61.9124,
  74.96166, 73.18517, 71.7793, 71.90649, 71.57249, 69.20923, 65.92067, 
    61.25922, 59.21616, 57.69858, 56.1347, 56.36287, 61.12395, 62.91213, 
    62.74499, 62.86666, 62.9311, 63.4561, 65.01925, 67.76344,
  94.24854, 94.52619, 94.71021, 94.95428, 94.98252, 95.0041, 95.37112, 
    95.47198, 94.23904, 94.40784, 94.3096, 94.30553, 94.40968, 94.28279, 
    94.44395, 94.96408, 93.79296, 93.82479, 93.82325, 93.92695,
  90.87362, 91.56668, 92.3815, 92.7374, 93.34521, 93.99747, 94.4807, 
    94.96357, 91.23316, 91.8055, 92.53537, 93.01187, 93.43978, 93.92699, 
    94.3167, 94.81979, 92.8513, 93.22023, 93.45986, 93.78307,
  85.89754, 87.31728, 88.54906, 89.80263, 90.87113, 91.73344, 92.95167, 
    93.58636, 89.04638, 89.69793, 90.193, 90.72643, 91.2628, 91.95036, 
    92.70208, 93.47907, 91.68964, 92.16913, 92.65766, 93.20757,
  84.02364, 85.27372, 87.1759, 88.4404, 89.91096, 91.24532, 92.73431, 
    93.82423, 90.93354, 91.36941, 92.02979, 92.34222, 92.85859, 93.09435, 
    93.49451, 93.6701, 94.6017, 94.77383, 95.21223, 95.17145,
  82.79347, 85.0115, 86.72578, 88.47762, 90.0591, 91.62582, 92.91167, 
    93.89532, 92.54554, 93.01857, 93.65035, 94.31761, 94.66861, 95.07578, 
    95.19145, 94.99395, 98.87023, 98.78598, 98.50424, 97.70413,
  82.11063, 84.61525, 86.69898, 88.33219, 89.31007, 90.39085, 91.17799, 
    92.03918, 87.96297, 88.22791, 89.17525, 89.84013, 90.26662, 91.4178, 
    92.53281, 93.91299, 99.43096, 99.55769, 99.50053, 99.24126,
  90.49549, 87.20533, 86.57793, 87.29435, 87.46681, 87.19703, 86.89441, 
    86.68919, 78.66783, 77.72627, 75.64886, 77.73542, 78.94906, 82.60361, 
    85.10881, 87.81787, 95.57988, 97.82826, 98.93504, 99.34542,
  93.15614, 93.07027, 93.33878, 93.50098, 93.64911, 93.22201, 92.7542, 
    92.39735, 85.39204, 82.71421, 77.11837, 81.07288, 82.00716, 87.78983, 
    82.31299, 75.3373, 75.48201, 92.71635, 93.40524, 95.26853,
  88.47466, 87.65739, 87.45789, 87.59064, 87.46294, 87.36782, 87.28247, 
    87.15417, 84.08415, 84.50036, 84.45933, 83.85231, 84.40697, 86.63625, 
    89.61641, 90.81059, 90.66386, 88.61787, 90.95114, 94.06027,
  91.60278, 91.53734, 90.92137, 89.60126, 87.68066, 85.5567, 84.79621, 
    84.11356, 83.86297, 84.44208, 85.9774, 87.78851, 89.04404, 90.62584, 
    91.81409, 92.87376, 93.50993, 94.36442, 94.71748, 94.69748,
  92.80476, 93.12881, 93.00933, 92.38747, 90.98682, 88.74939, 86.72816, 
    85.26031, 84.15463, 83.2071, 83.29533, 83.92522, 84.9246, 85.40242, 
    85.26013, 83.94537, 83.74618, 85.31365, 87.47445, 90.45946,
  92.23891, 92.27498, 92.19693, 91.91018, 91.56037, 90.32678, 88.72218, 
    88.02608, 87.06941, 85.15586, 83.25708, 82.54043, 83.70637, 85.08839, 
    85.21263, 84.33049, 83.1348, 82.72233, 83.90688, 85.74084,
  89.76324, 89.80893, 90.06149, 90.31898, 90.1101, 88.74474, 86.41775, 
    85.98074, 86.0591, 84.66537, 81.16354, 78.74287, 79.2485, 81.97554, 
    83.40617, 85.02059, 86.69546, 87.42889, 87.37383, 86.90577,
  88.95473, 88.68917, 89.07236, 88.65324, 85.96667, 82.75322, 80.4037, 
    79.43357, 79.07125, 79.7159, 79.9023, 80.13271, 80.78197, 82.74546, 
    84.64973, 85.59793, 85.82819, 86.82659, 88.0783, 88.74231,
  87.42553, 87.52565, 87.32481, 85.87194, 82.27695, 79.24329, 77.40044, 
    76.6078, 76.64035, 78.32711, 80.2008, 81.89638, 83.68416, 85.11069, 
    85.59048, 85.46106, 84.59788, 84.38007, 85.77503, 88.55721,
  84.64345, 85.00053, 83.21649, 79.49889, 76.26669, 75.19886, 75.22581, 
    75.54204, 76.17397, 78.44191, 80.99913, 83.32808, 85.12241, 86.2307, 
    85.62996, 84.31086, 83.25465, 82.89393, 83.80781, 85.34551,
  80.17444, 78.92461, 76.35806, 73.65244, 72.81552, 73.87192, 75.08165, 
    75.81384, 76.44608, 78.15523, 80.28677, 82.39327, 84.04502, 84.85776, 
    84.44993, 83.23632, 81.13928, 79.13005, 77.63445, 77.10226,
  75.67785, 74.29699, 73.6983, 72.74062, 73.60109, 74.16605, 73.33994, 
    70.2991, 66.05166, 65.42301, 67.70975, 71.43742, 74.85683, 76.7903, 
    77.54639, 77.36935, 74.5408, 71.07737, 69.29963, 69.51548,
  73.97976, 74.12706, 73.5762, 72.34396, 72.81382, 71.60871, 67.75245, 
    62.77557, 58.45661, 56.40585, 57.30446, 60.54505, 64.519, 67.41328, 
    68.8276, 68.83526, 68.03854, 67.44611, 67.53806, 68.30674,
  73.23138, 72.8726, 70.92344, 69.93272, 70.24886, 68.81299, 65.79192, 
    59.9808, 60.19387, 60.75865, 61.65036, 62.7752, 68.84103, 71.85408, 
    71.16816, 70.42018, 70.03639, 69.96913, 70.10913, 70.49166,
  89.96052, 90.14127, 90.46198, 90.68712, 90.94214, 91.16507, 91.35203, 
    91.62174, 90.27164, 90.43895, 90.56673, 90.90753, 91.1312, 91.3621, 
    91.52261, 91.72457, 90.97654, 91.20711, 91.36886, 91.62387,
  87.50953, 88.27721, 89.06524, 89.98952, 90.75108, 91.40243, 92.00845, 
    92.65055, 89.13295, 89.71069, 90.3354, 90.85617, 91.36628, 91.85039, 
    92.22512, 92.63766, 90.6228, 91.09321, 91.61871, 92.09299,
  84.27772, 85.51655, 86.65889, 87.94914, 89.10548, 90.44812, 91.49924, 
    92.52869, 88.18035, 89.21223, 90.08566, 90.94499, 91.68355, 92.69724, 
    93.50169, 94.1787, 92.25836, 92.8278, 93.25378, 93.72539,
  82.46832, 83.5116, 84.62366, 85.53696, 86.43139, 87.30471, 88.33424, 
    89.79129, 87.51632, 88.41357, 88.68939, 89.40958, 90.3707, 91.39353, 
    92.16387, 92.85557, 94.35446, 94.6618, 94.64343, 94.31229,
  82.04571, 83.89734, 85.63048, 86.95171, 88.08214, 89.30428, 90.3501, 
    91.25134, 89.52647, 89.71177, 90.19984, 90.25189, 90.45007, 90.45784, 
    90.38853, 90.41341, 94.86158, 94.59816, 94.02409, 93.11935,
  81.31824, 83.73799, 85.82955, 87.37961, 88.40699, 89.19422, 89.79917, 
    90.59454, 86.91176, 87.28291, 88.02271, 88.85509, 89.50159, 90.08857, 
    91.1856, 92.19197, 97.88627, 98.11152, 98.1786, 97.90118,
  87.85007, 84.34698, 83.33893, 84.11695, 84.64178, 84.56559, 84.41793, 
    84.10776, 76.34631, 76.00782, 75.60174, 76.56557, 78.66698, 83.88521, 
    86.43086, 86.95521, 94.316, 96.5034, 97.71924, 97.74382,
  89.91373, 88.37077, 86.52997, 84.87637, 83.29778, 81.43448, 78.5467, 
    76.11584, 67.96156, 66.3705, 66.60194, 72.19604, 72.19496, 74.0659, 
    67.40295, 70.89642, 74.29356, 93.71909, 92.48576, 94.01751,
  82.80268, 80.6633, 78.29031, 77.41553, 77.33784, 77.67278, 77.86601, 
    78.32744, 77.11636, 78.64951, 80.42534, 83.12768, 85.37569, 86.27148, 
    86.4593, 87.427, 88.66905, 88.59448, 92.04562, 95.18604,
  83.62095, 81.27309, 78.90241, 76.7127, 75.86523, 75.6237, 76.24973, 
    78.40787, 81.66679, 83.9035, 86.00951, 88.19665, 90.27612, 91.41143, 
    91.95866, 92.50025, 93.15086, 93.05527, 92.65839, 92.0948,
  86.25041, 85.98586, 85.35361, 84.16412, 83.25988, 82.73538, 82.78568, 
    83.76433, 85.57321, 86.60501, 87.10822, 87.68942, 88.77863, 89.46657, 
    89.02607, 87.95509, 88.17065, 89.11079, 89.89477, 90.60143,
  87.98073, 87.31393, 87.31535, 88.51035, 89.32664, 89.13741, 88.90334, 
    89.32542, 89.73669, 89.18324, 88.12354, 87.68253, 88.68317, 90.0575, 
    91.10783, 91.20965, 91.31303, 91.16023, 91.14361, 90.9493,
  89.22861, 88.01035, 87.55623, 88.31245, 89.26414, 88.57328, 87.05277, 
    87.39772, 88.69629, 88.51105, 87.12411, 86.06967, 86.24462, 88.46109, 
    90.64644, 91.87325, 93.28851, 94.18188, 94.17434, 93.47668,
  90.12554, 89.29005, 89.08926, 88.46768, 85.90206, 82.70692, 80.35603, 
    80.06805, 81.6105, 83.32106, 84.29008, 85.35744, 86.35052, 87.9183, 
    90.50227, 91.86723, 92.17172, 92.65219, 93.63606, 94.10207,
  89.63902, 88.8769, 87.79586, 85.4295, 81.70535, 78.94439, 77.2048, 
    77.32159, 79.09764, 81.30327, 83.44225, 85.80714, 87.90128, 89.52529, 
    90.77798, 91.28622, 90.73477, 89.77023, 90.32009, 91.9734,
  86.83028, 86.19446, 83.67227, 79.70783, 76.19196, 74.66554, 74.71467, 
    76.11174, 78.70892, 81.57884, 84.48672, 87.23185, 89.243, 90.33833, 
    89.97455, 89.0417, 87.8479, 86.83016, 87.16628, 87.76904,
  83.23926, 80.88559, 77.26088, 74.20995, 73.01216, 73.50414, 75.01592, 
    76.74947, 78.43192, 80.07734, 82.32954, 84.83373, 86.27312, 86.90289, 
    86.34198, 85.19165, 82.86086, 80.62987, 79.20681, 78.96643,
  79.76794, 76.90556, 75.18951, 74.5896, 75.22292, 75.8473, 74.51369, 
    70.37807, 66.45824, 66.24029, 69.02874, 72.60129, 74.92946, 76.61938, 
    77.30122, 77.22362, 75.19358, 73.37234, 73.62406, 75.55257,
  76.96545, 76.01836, 75.6974, 75.26392, 74.19289, 71.22932, 66.46104, 
    61.45201, 58.86634, 58.58348, 59.12359, 61.07524, 64.56969, 68.44405, 
    71.56593, 73.20352, 73.94464, 74.96944, 77.16821, 79.03782,
  72.04165, 71.17809, 70.06575, 68.55375, 67.73075, 66.21436, 64.43908, 
    60.98404, 62.98931, 65.642, 65.89089, 66.03248, 70.28543, 74.32901, 
    75.85719, 76.95969, 77.94371, 78.40154, 78.90559, 79.24483,
  88.14669, 88.48545, 88.96019, 89.33949, 89.74594, 90.05877, 90.37841, 
    90.70551, 89.31861, 89.69756, 90.0636, 90.36817, 90.65975, 90.91029, 
    91.21101, 91.4265, 90.63638, 90.85951, 91.02003, 91.1832,
  85.62018, 86.71167, 87.68246, 88.90178, 90.08609, 91.00537, 92.00358, 
    92.85702, 89.54574, 90.35345, 91.13479, 91.85405, 92.47932, 93.31144, 
    94.02507, 94.70218, 92.83823, 93.4285, 93.79006, 94.44512,
  85.16523, 86.46397, 87.87104, 89.34739, 90.7841, 91.97473, 93.1861, 
    94.23708, 90.11086, 91.15041, 92.10706, 93.13167, 94.25641, 95.29844, 
    96.15238, 96.97352, 95.34346, 95.9003, 96.42488, 96.87111,
  85.82774, 87.50355, 89.14076, 90.41764, 91.90329, 92.86704, 93.78461, 
    94.70528, 92.36752, 93.27709, 94.12395, 95.3126, 96.34225, 96.97701, 
    97.33902, 97.5637, 98.33056, 98.15899, 97.68541, 97.44537,
  85.44559, 87.93214, 90.10148, 91.98863, 93.15577, 94.26082, 95.11369, 
    95.70413, 94.8139, 95.39147, 95.99667, 96.26256, 96.60878, 96.86948, 
    96.88243, 96.78617, 99.37106, 99.14707, 98.48038, 97.71167,
  84.31215, 87.17559, 89.45306, 90.92074, 92.0005, 92.68012, 93.23607, 
    93.26405, 88.92326, 89.16837, 89.50817, 90.13419, 91.27751, 92.49881, 
    93.56751, 94.48876, 99.06667, 98.91228, 98.57707, 97.98473,
  90.99564, 89.07006, 88.45377, 88.16931, 87.74505, 87.44138, 87.01045, 
    86.49606, 78.44234, 78.31232, 78.25455, 78.11661, 79.42593, 85.20704, 
    88.42274, 85.83923, 93.13389, 95.43108, 96.65283, 96.99934,
  78.82176, 74.96894, 71.2406, 68.27242, 67.45467, 67.68376, 68.28155, 
    67.97612, 61.92902, 60.92236, 60.84499, 64.88483, 65.12808, 72.71735, 
    73.54975, 75.962, 81.84809, 90.44759, 89.95307, 91.73154,
  75.35437, 72.40674, 69.952, 68.22353, 67.76482, 68.82192, 70.20786, 
    71.63118, 70.62575, 71.39799, 72.60544, 74.08585, 76.08832, 78.67867, 
    80.15758, 79.80821, 78.37489, 75.28189, 83.66866, 90.74086,
  81.45335, 78.81551, 76.02112, 74.69998, 74.77735, 75.56722, 76.37621, 
    77.56741, 79.4951, 80.39996, 80.85433, 81.59937, 81.7817, 82.049, 
    82.71417, 83.28373, 83.85678, 83.8238, 83.68837, 83.89876,
  85.38638, 84.8242, 83.8994, 83.16936, 82.3429, 82.71018, 83.88361, 
    84.33477, 84.72235, 84.37307, 84.11703, 84.45689, 85.04396, 85.31155, 
    85.44554, 84.92144, 84.23567, 84.70358, 86.03726, 86.76934,
  90.51166, 90.49232, 90.47507, 90.5178, 90.48993, 90.02252, 90.01105, 
    90.05753, 89.48114, 88.56638, 87.43192, 87.09474, 87.84515, 88.72366, 
    89.27927, 89.27175, 88.69088, 88.68324, 89.51574, 90.27601,
  92.09871, 91.85294, 91.68975, 91.93927, 92.17593, 90.95555, 89.53798, 
    89.68539, 90.59967, 90.54823, 89.31359, 87.97951, 87.33917, 88.20467, 
    89.67263, 90.21435, 90.66235, 90.91199, 91.0424, 91.29337,
  91.07706, 90.64649, 90.79782, 90.80378, 88.83839, 86.82595, 85.88888, 
    85.61587, 85.97195, 86.62527, 86.71686, 86.8529, 87.35528, 87.80786, 
    88.84492, 89.20114, 88.75848, 88.93855, 90.07253, 91.17497,
  89.19271, 89.2251, 89.10001, 88.14419, 85.77593, 84.15875, 83.19487, 
    82.73212, 82.91482, 84.22668, 85.78731, 87.43301, 88.94386, 89.44718, 
    89.15278, 88.79527, 87.82008, 87.1386, 88.00566, 89.79023,
  84.55888, 84.79762, 83.67177, 81.37319, 79.17282, 78.57055, 78.8787, 
    79.54375, 81.22945, 83.6981, 85.96201, 88.03026, 89.22765, 89.43667, 
    88.04538, 86.8417, 85.55944, 84.99568, 85.67657, 86.17769,
  76.99928, 76.25504, 74.45943, 72.88246, 72.73112, 73.85565, 74.86557, 
    76.23796, 78.09113, 79.65154, 81.55938, 83.69639, 84.80418, 85.14212, 
    84.46414, 83.74498, 82.41752, 80.51747, 78.68659, 77.73586,
  70.03619, 68.93536, 68.91634, 69.68197, 71.05621, 71.8208, 70.27171, 
    67.06808, 65.53095, 65.85099, 67.40244, 71.0393, 75.32453, 77.77444, 
    78.3199, 78.01771, 76.01354, 73.16465, 71.22289, 71.33855,
  67.46931, 67.33266, 66.94579, 66.49998, 68.07883, 67.92564, 65.82078, 
    63.75012, 63.83933, 64.39008, 64.56578, 65.72561, 68.29697, 69.75941, 
    70.24621, 70.52374, 70.50028, 70.58622, 71.03468, 71.657,
  65.75106, 64.11977, 61.95403, 62.69769, 65.98875, 67.77412, 68.63983, 
    66.38372, 68.98563, 70.92297, 69.64422, 68.76864, 71.67599, 72.80981, 
    72.37975, 72.07307, 72.26851, 72.86623, 72.43641, 71.37982,
  92.38352, 92.75616, 93.11274, 93.49316, 93.7834, 94.03912, 94.42445, 
    94.83383, 93.43524, 93.74868, 94.10173, 94.35372, 94.81055, 94.91156, 
    95.38735, 95.5433, 94.71727, 94.73394, 94.74556, 95.45781,
  87.41257, 88.53493, 89.62611, 90.82851, 91.99921, 93.10319, 94.11863, 
    95.18478, 91.90836, 92.72742, 93.30348, 93.86174, 94.53339, 95.11552, 
    95.61068, 95.88765, 93.97594, 94.55096, 95.1855, 95.94463,
  83.03886, 84.68111, 86.32301, 88.02151, 89.55813, 90.94234, 92.15462, 
    93.26977, 88.81235, 89.35734, 89.74881, 90.38974, 91.75878, 93.35812, 
    94.92561, 96.15624, 95.26902, 96.43159, 97.47932, 98.31669,
  81.70889, 83.91233, 85.83372, 87.66615, 89.0866, 90.64723, 91.91508, 
    92.95479, 90.47989, 91.28489, 92.47778, 94.01394, 95.84386, 96.9957, 
    97.70159, 98.15102, 98.55312, 98.70299, 98.7756, 98.79906,
  80.08299, 82.85296, 84.96873, 85.67709, 85.74266, 86.96398, 87.42468, 
    88.44121, 88.1033, 89.14774, 90.12839, 92.31212, 93.65237, 94.70187, 
    95.35311, 95.79868, 98.2798, 98.19969, 97.84156, 97.41725,
  82.71856, 85.27038, 86.93849, 87.98216, 88.2438, 88.08386, 88.06501, 
    88.27974, 83.89013, 84.20039, 84.83284, 85.56542, 86.07995, 86.61815, 
    87.75111, 88.40819, 93.88446, 93.672, 93.81461, 93.39597,
  89.74101, 88.6405, 89.02799, 88.09132, 87.65829, 88.22886, 87.83031, 
    87.53934, 79.26507, 78.34486, 78.8572, 75.58064, 78.01794, 84.14127, 
    87.77858, 84.18359, 89.72059, 91.52219, 92.18402, 91.95191,
  71.28174, 70.34228, 68.83807, 65.15601, 64.3986, 66.35894, 65.92152, 
    64.50328, 58.96696, 58.14463, 60.12547, 67.29533, 73.00519, 81.64, 
    86.4536, 87.84875, 90.97649, 90.45611, 87.0729, 86.48443,
  69.27081, 68.64507, 69.3152, 69.84066, 70.41453, 72.00488, 73.86483, 
    75.60445, 75.75632, 77.46687, 78.21422, 77.87268, 77.13432, 77.53004, 
    78.15671, 78.93894, 81.80763, 86.39882, 89.72143, 92.66418,
  73.64888, 72.88657, 73.79284, 75.80708, 77.11349, 78.01984, 78.93888, 
    80.3001, 82.66229, 84.39886, 85.73035, 86.46738, 87.00554, 87.04293, 
    85.93878, 84.5424, 83.39005, 82.16202, 81.32211, 80.95684,
  80.1805, 79.93742, 79.92391, 80.34721, 80.36714, 80.5902, 81.40339, 
    82.28679, 84.18272, 85.34344, 86.33051, 87.24485, 88.02411, 88.43073, 
    88.05431, 87.11201, 86.53044, 85.99376, 85.57691, 85.26236,
  86.89226, 85.91376, 84.92686, 84.53689, 84.49162, 84.74917, 85.42999, 
    86.4828, 87.53165, 87.47925, 86.58972, 86.43842, 87.35678, 88.77718, 
    89.39855, 89.61194, 89.47012, 88.81322, 88.34828, 87.69538,
  89.60146, 88.75137, 87.90298, 87.64807, 87.5509, 86.63369, 85.51865, 
    85.65332, 86.66976, 87.01742, 86.02093, 85.51134, 85.72977, 87.24161, 
    89.81989, 91.24299, 91.43797, 91.20613, 90.74868, 89.84963,
  90.03717, 89.64641, 89.21038, 88.04417, 85.93365, 83.72775, 82.18493, 
    81.96803, 83.09338, 84.32724, 84.97756, 86.0948, 87.64583, 89.12135, 
    90.59241, 91.08424, 90.77386, 90.97713, 91.59117, 91.80719,
  88.90662, 88.80827, 88.18336, 86.27363, 82.89561, 80.6974, 79.82826, 
    80.33894, 81.63285, 83.47533, 85.45838, 87.56506, 89.40242, 90.41737, 
    90.69865, 90.51979, 90.44187, 90.71358, 91.62766, 92.82437,
  85.59312, 85.10937, 82.94569, 79.28434, 76.23039, 75.92147, 76.8735, 
    78.78367, 81.19417, 83.90374, 86.59187, 88.47067, 89.54501, 89.92414, 
    89.67728, 89.63869, 89.4544, 89.48494, 90.56818, 91.1421,
  77.76151, 75.53986, 73.04045, 71.23824, 71.00456, 72.47688, 74.7646, 
    77.05657, 79.11072, 81.07539, 83.27781, 85.30793, 87.03256, 88.41373, 
    88.28986, 88.01839, 87.60336, 87.20534, 86.85556, 86.55418,
  69.46916, 67.46565, 67.82101, 69.20148, 70.52895, 71.59665, 70.02895, 
    66.28799, 63.94594, 64.69608, 68.78482, 75.07005, 80.67629, 83.37454, 
    84.57394, 84.90273, 83.91223, 81.37933, 78.86056, 77.29759,
  67.28982, 67.8235, 68.1291, 67.9075, 67.55901, 66.03916, 63.43545, 
    61.11232, 61.52189, 61.67722, 64.07571, 68.5888, 72.72997, 73.7298, 
    73.53082, 73.1824, 72.72416, 71.90984, 71.82619, 71.57922,
  65.78514, 64.75299, 63.05461, 63.20816, 64.8064, 65.37786, 66.86034, 
    65.59279, 67.70692, 69.23982, 67.43883, 68.17059, 72.48109, 74.70657, 
    74.10088, 72.67375, 71.50545, 71.52197, 71.77389, 70.79636,
  94.09666, 94.45692, 94.85088, 95.30399, 95.64883, 95.96222, 96.2903, 
    96.51229, 94.96735, 95.42207, 95.74036, 95.82308, 96.11742, 96.43303, 
    96.74052, 97.00308, 95.93322, 95.93768, 96.17094, 96.67374,
  88.94659, 90.0891, 91.18869, 92.14777, 93.19633, 93.88898, 94.70737, 
    95.38248, 92.0146, 92.68272, 93.36264, 93.95062, 95.00563, 95.51551, 
    96.21117, 96.35178, 94.79522, 95.2786, 95.92713, 96.46254,
  88.44798, 89.84161, 91.44447, 92.86613, 94.05758, 94.84141, 95.89102, 
    96.56462, 92.28883, 93.15574, 94.16216, 95.11598, 95.68926, 96.2826, 
    96.3549, 95.9556, 94.74216, 95.33549, 96.3086, 97.21377,
  86.73839, 88.87447, 90.96143, 93.2722, 95.30807, 96.59537, 97.75264, 
    98.49114, 97.16405, 97.84389, 98.48356, 98.68918, 98.19562, 98.46701, 
    99.22945, 99.66016, 99.80584, 99.8621, 99.77495, 99.22205,
  80.9132, 83.22937, 85.21889, 87.46844, 89.74955, 90.8001, 92.52611, 
    93.76968, 93.5309, 94.3895, 94.71523, 94.78459, 95.72762, 96.66558, 
    97.46224, 98.22386, 99.66812, 99.83062, 99.7823, 99.74133,
  81.00658, 83.76553, 85.60507, 86.15141, 87.15131, 87.35083, 87.29234, 
    86.73335, 82.15459, 82.36114, 82.95345, 84.0141, 85.52016, 86.92798, 
    88.05162, 88.75213, 95.19517, 96.29781, 97.07104, 96.95768,
  93.7969, 89.54942, 89.75323, 90.26025, 90.22526, 89.84125, 89.02749, 
    87.94978, 79.72536, 79.98832, 81.31232, 77.28825, 78.21809, 81.48618, 
    86.27432, 81.48704, 87.19439, 89.65228, 91.76204, 93.14305,
  76.29688, 76.06165, 77.28992, 79.33677, 80.81233, 82.74747, 83.32902, 
    82.9877, 75.38077, 75.55396, 77.78858, 74.78378, 77.19102, 83.38418, 
    91.27814, 91.19852, 93.16972, 91.19785, 90.17165, 89.88238,
  68.08606, 65.47161, 63.37497, 62.14815, 62.0598, 62.5656, 62.62481, 
    62.23506, 59.24091, 61.25058, 65.24506, 72.28333, 79.16814, 82.77416, 
    84.04621, 85.15948, 88.17433, 91.38102, 93.27881, 93.76263,
  75.60804, 73.56903, 71.64053, 69.57486, 68.3282, 67.41896, 66.81322, 
    66.0048, 64.96113, 64.68983, 65.12505, 66.31941, 67.78487, 69.46472, 
    71.17119, 73.24031, 76.39331, 78.5292, 79.62492, 80.19534,
  82.42992, 81.1775, 79.43147, 76.90778, 74.50888, 73.14402, 72.63885, 
    72.35605, 71.80772, 71.34604, 71.35997, 71.98389, 73.07014, 74.10029, 
    74.71455, 75.46703, 77.32571, 78.53448, 79.25942, 80.29972,
  86.82232, 86.36077, 85.18151, 83.29557, 81.29726, 79.53965, 78.41044, 
    77.85994, 76.84786, 75.42757, 73.71926, 73.22776, 74.29282, 76.08884, 
    77.46995, 78.0743, 79.01866, 79.96177, 81.13455, 82.29486,
  88.6201, 87.7767, 87.13017, 86.13629, 84.52139, 82.01437, 79.58067, 
    78.2564, 76.98048, 75.52438, 73.46303, 72.3019, 72.54823, 74.31515, 
    77.41405, 79.47314, 80.06659, 80.85662, 81.64453, 82.09872,
  88.76805, 88.37066, 87.75253, 86.07688, 83.43633, 80.67395, 78.11433, 
    76.23569, 74.76276, 74.04897, 73.18466, 72.78452, 73.42491, 75.32731, 
    77.85146, 78.87007, 78.0696, 78.1678, 79.61063, 80.89668,
  87.33857, 87.35947, 86.7523, 84.68212, 81.16548, 78.5361, 76.27422, 
    74.49054, 73.67097, 74.04359, 74.5551, 75.3952, 76.66356, 78.04336, 
    79.06286, 78.92274, 77.74725, 77.529, 78.87756, 81.31972,
  84.14855, 84.36045, 82.64075, 79.28075, 75.8691, 74.59415, 73.96675, 
    73.86633, 74.28429, 75.90878, 77.70168, 79.08623, 80.05009, 80.6655, 
    80.25718, 79.57137, 78.42931, 77.78754, 78.71459, 79.98426,
  77.64831, 76.3028, 73.79535, 71.21865, 70.71024, 72.48446, 74.85023, 
    76.44572, 77.20466, 78.21602, 79.52008, 80.61777, 81.26102, 81.26743, 
    80.52642, 79.41593, 77.38378, 75.70861, 75.05434, 75.55887,
  69.1367, 66.77879, 68.00219, 70.27119, 72.67355, 74.50442, 72.8447, 
    68.11952, 65.76066, 66.07876, 68.21827, 71.14182, 73.42954, 73.86694, 
    73.85461, 73.65705, 71.62498, 69.7794, 69.89555, 71.45174,
  65.27884, 66.79971, 69.52439, 71.52027, 71.75895, 68.66898, 64.96552, 
    63.20227, 62.79242, 60.80029, 61.14416, 62.40417, 63.62528, 63.31229, 
    62.81896, 63.51891, 64.76029, 66.09676, 68.10908, 70.58105,
  65.40778, 66.62852, 67.21, 67.79871, 68.37026, 68.53746, 68.7126, 65.36804, 
    64.66512, 63.99017, 61.516, 61.42529, 64.05882, 66.13109, 66.47616, 
    67.5342, 69.2951, 70.88873, 72.00098, 72.89951,
  91.83164, 92.12141, 92.38763, 92.63519, 93.07784, 93.29901, 93.59207, 
    93.95804, 92.59431, 92.95277, 93.42178, 93.74726, 94.16886, 94.21516, 
    94.768, 95.26431, 94.59103, 94.8558, 95.24256, 95.51273,
  86.98829, 88.03703, 88.85042, 89.70961, 90.99543, 92.27769, 93.53139, 
    94.4806, 91.6512, 92.6357, 93.66724, 94.47924, 95.23271, 95.52451, 
    95.77048, 96.12059, 94.41225, 94.88375, 95.52407, 96.31084,
  86.12935, 87.88772, 89.03889, 90.45998, 91.79535, 92.55376, 93.81791, 
    95.00117, 90.44573, 91.234, 92.47, 93.78156, 95.00211, 96.5443, 97.49848, 
    98.33726, 97.50896, 97.79507, 97.67779, 97.51231,
  85.98232, 88.86978, 91.15259, 92.71851, 93.40595, 94.05857, 94.72604, 
    95.1313, 92.68478, 93.26325, 94.04541, 95.1757, 96.39442, 97.75491, 
    98.80005, 99.08231, 99.36423, 99.49146, 99.57432, 99.53441,
  83.11666, 86.05652, 88.27755, 88.88128, 89.18862, 89.70999, 90.39392, 
    91.18778, 90.67983, 91.44788, 92.60716, 94.14944, 95.71284, 96.91077, 
    97.68313, 98.26732, 99.41599, 99.37527, 99.11376, 98.81631,
  84.96561, 87.31104, 88.60865, 89.02235, 89.05251, 88.7813, 88.83686, 
    88.77896, 84.52093, 84.63795, 84.95767, 85.83539, 86.46108, 86.88548, 
    87.16647, 88.51086, 95.84919, 96.74643, 97.36395, 97.17663,
  98.12476, 94.58668, 93.37181, 92.69833, 92.21141, 92.40253, 92.26414, 
    92.12928, 84.18534, 84.44837, 85.88981, 79.19331, 79.69906, 84.17367, 
    88.51752, 84.10229, 88.75932, 90.56798, 92.16796, 92.96539,
  98.66299, 98.05103, 96.14562, 93.10862, 92.75006, 94.06523, 94.60263, 
    94.31251, 89.99966, 89.90438, 90.89071, 86.13617, 86.80898, 90.32935, 
    95.20692, 93.92852, 94.81634, 93.00977, 91.11938, 92.1892,
  85.89071, 85.8866, 87.60736, 90.82909, 93.02747, 93.81869, 94.22981, 
    94.31105, 93.16946, 93.14752, 94.03171, 93.52833, 93.12781, 92.78002, 
    92.3571, 90.58652, 92.62516, 95.41046, 96.57793, 95.79547,
  72.90121, 75.80883, 78.5319, 79.85968, 81.38158, 83.55543, 84.21901, 
    83.78107, 82.50922, 81.17213, 80.39815, 78.88828, 76.27506, 73.45739, 
    71.73899, 73.02396, 77.0906, 82.53683, 88.08357, 89.08697,
  64.94266, 66.03613, 67.06956, 67.33932, 67.91877, 68.50288, 69.33553, 
    70.41994, 70.05769, 69.21371, 68.08162, 66.69553, 67.39079, 69.41706, 
    71.31425, 71.2019, 70.6244, 70.16872, 69.66235, 68.68525,
  58.83146, 59.00249, 59.18668, 60.37679, 62.12365, 63.84061, 65.05106, 
    66.89551, 68.51658, 68.98565, 68.57424, 68.84597, 70.63029, 74.06994, 
    77.14213, 78.19746, 77.80698, 76.84808, 76.0065, 74.8399,
  63.72718, 64.24766, 65.10673, 66.65717, 67.8166, 68.32167, 68.39661, 
    69.44736, 70.94319, 70.97652, 69.96781, 69.32037, 70.00298, 72.76164, 
    77.35158, 80.4146, 81.28554, 81.17341, 80.3928, 78.80566,
  72.29696, 71.85582, 71.89413, 71.40272, 69.46234, 67.45251, 66.39599, 
    66.55785, 68.20605, 69.55065, 69.72939, 69.98376, 71.13543, 73.8335, 
    77.33353, 79.70101, 80.23911, 80.1684, 80.50157, 81.28492,
  77.44198, 77.47758, 77.00235, 75.32017, 72.06982, 69.44899, 67.95972, 
    67.68742, 69.51147, 71.795, 73.7746, 75.51082, 77.18294, 78.87365, 
    80.44438, 81.32347, 80.97424, 80.14672, 80.713, 82.67675,
  77.43478, 77.70647, 76.11465, 72.45267, 68.86536, 67.24125, 67.32954, 
    68.67979, 71.61855, 75.00645, 78.53885, 81.48939, 83.66759, 84.9875, 
    84.58888, 83.2218, 81.62186, 80.93445, 81.92763, 83.18555,
  73.86352, 72.19901, 68.58063, 64.9032, 63.46404, 64.67788, 67.13621, 
    69.9874, 73.35418, 76.15806, 79.3171, 82.12319, 84.38319, 84.96326, 
    84.0368, 83.06799, 81.81458, 80.53932, 79.7366, 78.84282,
  66.97176, 64.26828, 64.63072, 66.71768, 68.66816, 70.34808, 68.52786, 
    63.58456, 60.54251, 60.94458, 64.13258, 69.20032, 74.04996, 76.6747, 
    78.14954, 78.8148, 77.23967, 74.54665, 72.82187, 71.88029,
  65.25487, 66.85786, 69.17866, 71.1076, 69.73647, 64.64542, 59.29459, 
    56.3503, 55.96213, 54.65669, 55.01846, 57.26001, 60.6534, 64.46171, 
    67.19821, 68.83735, 70.02711, 70.7583, 71.88963, 73.44189,
  67.46601, 67.52341, 67.29771, 66.07036, 63.84837, 62.04328, 61.08063, 
    61.84337, 62.06443, 61.05221, 56.53541, 57.12112, 62.15476, 67.23957, 
    69.72263, 71.03848, 73.13203, 75.68156, 78.3026, 79.57047,
  93.75117, 94.07439, 94.52319, 94.83181, 95.16676, 95.56477, 95.94667, 
    96.19295, 94.77646, 95.12841, 95.50146, 95.70948, 95.90677, 96.17332, 
    96.47986, 96.70333, 95.72953, 95.79858, 95.85405, 96.10705,
  90.21169, 91.05286, 91.93307, 92.71626, 93.5771, 94.16097, 94.94704, 
    95.47473, 92.01492, 92.46819, 92.94088, 93.59775, 94.09661, 94.62048, 
    94.60368, 95.59811, 93.7563, 95.8595, 96.60905, 97.39289,
  88.76234, 90.19202, 91.63408, 93.01128, 94.63845, 95.30228, 95.89523, 
    96.47669, 92.05225, 92.92103, 93.66935, 94.87624, 96.19638, 97.30701, 
    97.81854, 98.40285, 97.81538, 98.15678, 98.36341, 98.68151,
  87.29491, 89.55466, 91.354, 92.98414, 94.38271, 95.53609, 96.9904, 
    97.93634, 95.80942, 95.9571, 96.04626, 96.33118, 96.83769, 97.56098, 
    98.42725, 98.76237, 99.13856, 99.29913, 99.1655, 98.617,
  87.42381, 89.85838, 91.78887, 93.01543, 93.81588, 93.81563, 94.08246, 
    94.53569, 94.09802, 94.66076, 95.59034, 96.41481, 97.06409, 97.53161, 
    97.62348, 97.48525, 98.94334, 98.98624, 99.11316, 99.13802,
  82.69518, 85.08162, 86.81229, 87.57292, 87.21968, 87.4363, 87.84623, 
    88.27322, 84.50474, 84.6804, 84.19138, 84.84417, 86.306, 88.05423, 
    89.93761, 91.73595, 97.63239, 98.34814, 98.8166, 98.69856,
  94.44095, 87.73863, 86.81301, 87.40799, 87.19794, 87.25136, 87.67357, 
    87.99297, 80.35573, 80.47158, 82.13231, 77.81148, 79.18409, 84.5008, 
    87.57627, 86.38206, 92.34182, 94.2452, 95.22163, 95.582,
  96.47829, 96.36175, 97.28665, 97.74479, 97.14309, 96.96764, 96.19781, 
    95.77322, 92.08547, 92.29411, 94.19829, 89.77232, 89.6715, 92.38863, 
    94.70197, 93.67336, 94.60599, 95.80363, 92.99068, 94.73027,
  96.0071, 96.04324, 95.7799, 95.25349, 95.65176, 95.48456, 95.54796, 
    95.88134, 95.93301, 96.89312, 97.26216, 97.25372, 96.60629, 95.8389, 
    96.08998, 96.17414, 97.12549, 98.14745, 98.57537, 98.91258,
  95.45307, 94.35132, 94.89982, 95.6735, 95.76952, 95.90862, 95.72151, 
    96.06433, 96.3133, 96.87176, 96.60635, 96.07948, 95.36794, 95.45313, 
    94.75361, 93.51543, 93.89716, 95.58736, 97.0218, 97.98225,
  94.4063, 94.48646, 95.15366, 95.63236, 96.18428, 96.35405, 96.6926, 
    96.32272, 95.30666, 92.98053, 91.15077, 89.89931, 86.02715, 82.21122, 
    79.59899, 76.75465, 74.81129, 75.27605, 77.86337, 79.16875,
  85.40729, 85.98556, 86.40366, 87.79143, 87.51572, 86.02858, 82.7355, 
    78.49966, 71.88865, 66.97613, 64.52254, 63.90934, 64.48989, 66.47938, 
    68.70012, 69.61585, 69.91245, 70.38432, 70.53838, 69.97697,
  64.29028, 64.12489, 65.11015, 66.89439, 68.06496, 68.45723, 67.99889, 
    68.07061, 68.36626, 68.1171, 67.37793, 66.98877, 66.85231, 67.85246, 
    70.46468, 73.36236, 75.04635, 76.35783, 77.16435, 76.63099,
  67.48267, 67.84632, 68.83635, 69.20768, 68.36809, 67.45683, 67.08226, 
    67.39543, 68.5142, 69.62772, 70.29002, 71.03929, 72.09701, 73.85453, 
    76.82346, 79.62165, 80.88974, 81.94081, 83.08088, 83.20071,
  70.03927, 70.79227, 71.24141, 70.38334, 68.22485, 66.58235, 65.24632, 
    64.70566, 66.15609, 68.56885, 71.28541, 74.60526, 77.63826, 80.18301, 
    82.76964, 84.4882, 84.7346, 84.19713, 84.59737, 85.59721,
  69.45535, 70.49178, 69.5839, 66.83484, 63.58308, 61.83027, 61.27952, 
    62.15477, 65.69614, 70.49722, 75.2973, 79.59803, 83.26157, 85.79988, 
    86.6242, 86.38812, 85.22056, 83.98437, 84.28196, 84.8268,
  66.28166, 64.57861, 61.84436, 58.90305, 56.85143, 57.66194, 60.12186, 
    63.5202, 68.12835, 73.00928, 78.06289, 82.29424, 85.35522, 86.88717, 
    86.38107, 85.57814, 83.83086, 81.75935, 80.08934, 78.84508,
  58.14913, 55.00607, 54.91447, 56.90548, 59.85913, 63.27074, 64.71404, 
    62.80013, 61.92972, 63.47636, 67.21457, 71.63913, 75.62054, 78.16718, 
    79.02945, 79.10426, 76.81431, 72.71773, 69.93169, 69.20176,
  60.16754, 61.76697, 64.13488, 66.61622, 67.21008, 63.7873, 59.23803, 
    56.97776, 57.36765, 56.13837, 56.81221, 59.21848, 62.92901, 65.68423, 
    67.00322, 66.62217, 65.68425, 63.95539, 63.54333, 64.70094,
  69.09082, 70.10526, 69.91185, 68.50211, 65.36502, 62.33908, 61.51354, 
    61.31862, 62.59515, 61.0095, 57.24099, 58.30297, 64.66415, 69.23987, 
    70.18071, 69.16703, 68.4564, 67.9221, 69.30932, 71.43628,
  91.63286, 92.06338, 92.2374, 92.90601, 93.22282, 93.57597, 94.13648, 
    94.75221, 93.1732, 93.44183, 93.66608, 94.30631, 94.74939, 94.97086, 
    95.24662, 95.68503, 94.58875, 94.63612, 95.2999, 95.26384,
  85.36668, 86.79665, 88.28246, 89.91779, 91.42029, 92.98025, 94.0276, 
    95.23365, 91.48306, 92.49756, 93.19638, 94.01501, 94.54793, 95.64721, 
    95.91011, 97.62363, 96.55145, 97.29047, 97.54023, 97.99926,
  84.31036, 86.17881, 88.19482, 90.13496, 91.56853, 92.8563, 93.83437, 
    95.12043, 90.5895, 92.46429, 93.79667, 95.1461, 96.17406, 97.15369, 
    98.23701, 98.68761, 98.23164, 98.09296, 97.82457, 98.16542,
  85.29055, 87.67006, 90.13828, 93.15862, 95.00861, 95.83928, 96.1486, 
    96.16268, 94.0228, 94.468, 95.95217, 97.1382, 97.74272, 98.14603, 
    98.5223, 98.93166, 99.34424, 99.30342, 98.97874, 99.01895,
  83.83271, 86.41897, 88.3604, 89.43664, 90.39893, 91.52729, 91.81873, 
    91.58489, 91.26922, 92.02098, 93.0399, 93.58141, 94.01893, 94.35016, 
    95.59361, 96.44323, 98.81899, 98.50191, 98.32179, 98.16138,
  79.48873, 82.06803, 84.76179, 87.35992, 89.5363, 91.10649, 92.44963, 
    92.60262, 86.3724, 86.02383, 86.40332, 88.07306, 89.72739, 91.18056, 
    92.62164, 94.04927, 98.87597, 98.98737, 98.32246, 96.79226,
  98.08701, 92.82185, 93.67473, 93.96488, 93.14211, 92.62981, 91.73292, 
    91.1188, 83.20451, 83.75301, 85.32292, 79.12861, 81.14196, 88.95309, 
    91.41604, 88.6992, 94.45396, 94.54344, 94.68024, 93.77622,
  97.45689, 97.55807, 97.38981, 97.10332, 97.23473, 97.32471, 97.23351, 
    97.12206, 95.00217, 95.26892, 96.62238, 93.82697, 93.79216, 96.3347, 
    97.87494, 91.438, 97.06296, 97.24776, 93.86063, 94.60281,
  97.36477, 97.52534, 97.42724, 97.88829, 97.99876, 98.3226, 98.66637, 
    98.00581, 95.7903, 96.43265, 97.88769, 99.47272, 99.33215, 99.05059, 
    98.46079, 98.37109, 98.53651, 99.37896, 99.44541, 98.33414,
  96.25, 96.59024, 97.37301, 97.50086, 97.12793, 96.53779, 95.73576, 
    94.78792, 93.79902, 93.14561, 94.93325, 97.27878, 97.79958, 97.62624, 
    97.18201, 97.3671, 97.64046, 98.24799, 98.63467, 98.63454,
  95.57013, 97.30104, 97.72841, 97.86516, 97.83369, 97.76589, 97.03439, 
    96.01001, 96.13023, 96.31955, 96.01865, 95.3257, 94.73259, 94.50165, 
    94.10139, 94.40943, 93.7554, 93.68116, 94.4689, 95.18658,
  95.36193, 96.12533, 96.54244, 97.04773, 97.0699, 96.32604, 95.91867, 
    95.17421, 93.91627, 80.64725, 67.47743, 62.4346, 62.45994, 66.09969, 
    69.8842, 78.68372, 86.30095, 89.05676, 87.17725, 85.19568,
  87.58375, 85.27862, 85.45441, 82.84837, 77.85686, 72.27901, 66.58263, 
    63.99475, 62.75067, 59.52407, 57.49512, 56.86342, 57.15872, 58.40632, 
    61.01309, 63.73408, 66.48619, 68.50566, 69.82958, 68.58379,
  67.82051, 66.81849, 66.26481, 64.62408, 62.41994, 60.4606, 58.49615, 
    57.49258, 57.93657, 59.34562, 60.01577, 60.59943, 62.16097, 64.28761, 
    66.94769, 69.38842, 70.23147, 71.06614, 72.28614, 73.36877,
  70.20546, 69.21955, 67.94164, 65.72917, 62.52405, 59.80277, 57.02002, 
    55.14744, 55.15827, 57.06247, 59.93415, 63.24844, 66.70243, 69.58163, 
    71.92043, 73.7323, 74.54377, 74.93545, 76.44479, 78.64719,
  73.55582, 71.92899, 68.62239, 64.02635, 59.92204, 57.57882, 55.59732, 
    54.3631, 55.48772, 59.28011, 64.75887, 69.93781, 73.46526, 76.26795, 
    78.65594, 79.59299, 79.15062, 78.32817, 78.95131, 80.27612,
  71.29507, 67.19216, 61.57364, 57.08992, 55.34027, 55.37474, 56.20221, 
    57.70671, 60.54174, 65.2104, 70.27213, 74.17278, 77.50191, 80.078, 
    81.59105, 81.79813, 80.44764, 78.47514, 76.78173, 75.71436,
  62.07628, 57.638, 56.13784, 57.01241, 59.19507, 61.89791, 63.40826, 
    61.65807, 59.94757, 60.34737, 62.43775, 65.84382, 70.22263, 74.14484, 
    76.98451, 77.11186, 74.71877, 70.87019, 67.47521, 65.66759,
  62.71289, 63.47077, 65.47664, 68.31433, 69.40111, 66.51028, 61.65962, 
    58.9253, 57.3884, 54.3226, 53.59658, 55.4603, 59.33649, 63.14934, 
    65.23686, 65.44052, 64.31004, 62.52524, 61.88379, 62.24872,
  72.066, 72.29118, 72.09295, 70.82845, 66.84677, 62.52596, 60.99018, 
    61.49741, 61.04218, 58.15757, 52.80347, 53.61164, 60.5975, 65.99304, 
    66.87312, 66.51982, 66.44012, 66.73515, 67.90155, 69.00552,
  93.3803, 93.78398, 94.16505, 94.41261, 94.55999, 94.95307, 95.15911, 
    95.44941, 93.97588, 94.37879, 94.58595, 94.85509, 95.1852, 95.40089, 
    95.71676, 96.05057, 95.32906, 95.43505, 95.51796, 95.66494,
  89.2565, 90.39099, 91.47807, 92.54034, 93.40849, 94.11253, 94.92072, 
    95.68069, 91.93992, 92.72108, 93.51672, 94.40727, 95.32605, 96.02582, 
    96.58257, 97.12115, 95.98985, 96.81357, 97.42504, 97.81281,
  89.94517, 91.01814, 91.91574, 92.7121, 93.36819, 94.15925, 94.7066, 
    95.32845, 90.42682, 91.34406, 93.37688, 94.58215, 95.12056, 95.95266, 
    96.07108, 96.34402, 96.09533, 97.34756, 98.06606, 98.55437,
  87.97871, 89.48976, 91.2726, 92.89738, 93.67667, 94.8335, 95.65894, 
    96.58752, 95.01093, 95.15829, 94.66502, 94.92572, 96.01639, 98.66838, 
    99.37988, 99.55767, 99.54009, 99.38808, 99.37008, 99.38717,
  86.94555, 89.03905, 90.57217, 91.36924, 90.86996, 91.01746, 90.50639, 
    89.22938, 88.55936, 90.03949, 91.1838, 92.47062, 94.30068, 96.28029, 
    97.57334, 98.14597, 99.49799, 99.80679, 99.90231, 99.75073,
  86.72569, 87.80264, 87.77773, 86.13857, 85.18392, 85.03796, 85.61762, 
    87.07594, 83.85263, 85.17307, 86.70908, 88.42869, 90.05549, 91.76234, 
    93.27892, 94.36424, 98.68432, 98.99652, 99.16464, 99.41335,
  94.75902, 93.35898, 92.46275, 90.2988, 88.05312, 86.91174, 86.21673, 
    86.52379, 79.44021, 80.5679, 82.84807, 75.82074, 77.76267, 86.08567, 
    87.62339, 84.71941, 92.72318, 95.04967, 95.86222, 95.59811,
  99.31831, 98.98946, 98.55882, 98.12373, 96.77994, 95.86936, 96.31283, 
    97.14888, 92.68259, 93.65385, 94.39069, 93.8366, 94.90681, 97.89284, 
    97.9581, 90.38847, 96.57664, 97.08214, 91.53742, 92.70068,
  98.97001, 99.11275, 98.71693, 98.38494, 98.32878, 97.36066, 96.34287, 
    95.78233, 94.04199, 95.31451, 95.97033, 96.46999, 97.61996, 97.92735, 
    97.92408, 97.81915, 97.90266, 98.36436, 98.36639, 97.78177,
  96.76794, 96.90106, 96.90757, 96.8362, 96.86684, 96.80616, 96.50841, 
    96.74809, 97.09911, 97.27125, 97.27676, 97.32491, 97.21236, 97.38557, 
    97.75956, 97.51801, 97.29677, 97.10817, 97.12774, 97.15923,
  95.63883, 95.48675, 94.94024, 94.69298, 95.03556, 95.12946, 95.15281, 
    95.64554, 96.00769, 96.13791, 95.81339, 95.24223, 94.90782, 95.03806, 
    95.7084, 96.45539, 96.93163, 97.08386, 96.64541, 96.44168,
  95.0427, 94.96944, 94.7542, 94.68897, 94.66216, 94.6649, 94.21351, 
    93.67982, 92.71754, 91.39075, 86.4491, 80.50067, 77.08253, 78.62228, 
    87.17997, 91.2197, 93.22939, 94.36735, 94.40575, 95.25279,
  93.08722, 92.90386, 92.4191, 91.74494, 90.70801, 89.03935, 85.79826, 
    82.16906, 78.42256, 73.17454, 66.20958, 61.53675, 60.73081, 62.48849, 
    66.6332, 70.21813, 72.91339, 76.3334, 80.6357, 79.71461,
  85.78922, 84.44907, 82.56175, 79.21632, 75.1896, 71.44221, 68.63203, 
    67.17915, 66.2775, 66.05505, 64.88577, 64.32765, 65.81403, 68.25632, 
    70.48204, 71.88429, 71.69178, 71.89919, 72.55126, 72.96185,
  82.93491, 81.87, 79.80025, 76.38248, 71.61803, 68.39849, 66.33471, 
    65.04961, 64.68125, 65.73312, 67.08556, 69.23476, 71.97247, 73.70345, 
    74.1369, 74.58145, 74.81882, 74.61943, 75.03643, 76.10391,
  80.31142, 79.45883, 76.19868, 70.36041, 64.56038, 62.09403, 61.94048, 
    62.2217, 63.78482, 66.80492, 70.47066, 73.9538, 76.30766, 77.38846, 
    77.52903, 77.35442, 76.45647, 75.36044, 75.87109, 77.0912,
  74.58528, 70.51932, 64.79327, 59.58315, 56.79563, 56.79262, 57.91712, 
    59.53658, 62.1267, 65.60511, 69.50528, 73.17189, 75.80943, 77.83872, 
    78.70288, 78.15131, 76.1302, 74.15353, 72.80168, 72.12557,
  62.68829, 58.02236, 56.46438, 56.6259, 57.45908, 58.97396, 60.09055, 
    59.09647, 57.53768, 57.43649, 58.49759, 61.11096, 64.45536, 67.48717, 
    70.49821, 71.63092, 69.18011, 65.75128, 63.49504, 62.92969,
  57.47611, 59.12222, 61.32402, 63.34715, 64.38023, 62.97862, 59.57952, 
    57.28402, 55.78019, 53.67193, 52.53043, 53.32402, 55.52057, 57.77143, 
    59.82248, 61.03461, 60.7352, 59.76455, 59.50418, 60.17618,
  62.00339, 64.14494, 66.22587, 67.0239, 63.74706, 60.23272, 59.7207, 
    63.51487, 64.11444, 61.31556, 53.96448, 53.44645, 59.3903, 63.34978, 
    64.42979, 64.04398, 63.43678, 63.00071, 62.98062, 63.61975,
  91.36868, 91.90617, 92.46822, 92.76107, 93.26398, 93.69603, 94.12927, 
    94.5331, 93.36361, 93.88871, 94.32327, 94.62672, 95.01989, 95.01487, 
    95.67235, 96.10377, 95.63415, 95.7835, 95.82011, 96.01574,
  84.36562, 85.88667, 87.44104, 88.88521, 90.15939, 91.44559, 92.7226, 
    94.11312, 90.817, 92.07552, 93.21806, 94.09611, 95.28117, 96.49084, 
    97.47681, 98.5017, 97.91014, 98.59665, 99.1389, 99.50607,
  83.11755, 85.20869, 87.04724, 88.59719, 90.0796, 90.98827, 91.82798, 
    92.52222, 87.89717, 88.3725, 90.11216, 91.4147, 93.31327, 95.01175, 
    95.90166, 96.53723, 95.84597, 96.4108, 96.80576, 97.39907,
  79.04953, 81.10337, 82.87112, 84.92475, 86.70061, 87.4167, 88.31401, 
    89.20628, 87.58594, 89.39535, 91.67931, 94.28828, 96.1421, 97.04437, 
    97.56631, 97.73659, 97.87071, 97.5856, 97.34927, 96.9258,
  74.92532, 76.97306, 78.77195, 80.66471, 82.00155, 83.64912, 84.51775, 
    86.39679, 87.04541, 88.88669, 90.90873, 92.75442, 94.66763, 96.35024, 
    96.78641, 96.68053, 98.65122, 98.67822, 98.46206, 98.10232,
  75.68324, 77.51283, 79.03325, 79.66767, 80.88632, 82.06963, 83.26398, 
    84.24973, 80.58392, 81.45998, 82.80411, 84.49011, 86.44592, 88.43831, 
    90.04351, 91.4331, 96.77888, 97.32321, 97.64467, 97.47621,
  92.69888, 88.21475, 85.71321, 83.23145, 82.8077, 83.69064, 84.06484, 
    84.66368, 76.96703, 77.36066, 79.15868, 73.00421, 75.68867, 84.28, 
    85.33775, 85.00843, 92.28845, 93.99982, 95.307, 95.92377,
  97.44506, 97.08164, 95.80946, 93.8019, 95.14804, 96.50967, 97.02918, 
    97.7078, 92.95973, 93.15878, 95.78011, 94.68349, 95.33231, 97.39194, 
    98.5479, 88.71239, 96.74498, 94.76339, 93.51092, 93.91853,
  96.51432, 96.51257, 95.88793, 95.14474, 95.05869, 94.83281, 93.7506, 
    93.04797, 91.97343, 93.06179, 94.46175, 96.65237, 97.494, 97.70905, 
    98.16171, 98.46863, 98.58081, 99.07729, 98.99775, 98.69911,
  96.53839, 96.00578, 95.95117, 95.86388, 96.08764, 96.17911, 95.34766, 
    94.40314, 94.3972, 94.99283, 95.90039, 96.19324, 96.12991, 96.2653, 
    96.72377, 97.61919, 97.9245, 98.11723, 98.26722, 97.84292,
  96.55254, 96.49165, 96.55133, 96.42452, 96.14478, 95.99911, 95.32106, 
    94.95123, 95.5209, 95.79725, 95.57587, 95.0104, 93.91077, 93.57323, 
    93.90371, 94.5909, 94.31209, 94.58627, 95.88288, 96.49377,
  95.36266, 95.63879, 95.77309, 95.25513, 94.76192, 94.24618, 94.14989, 
    94.24942, 93.95879, 94.13154, 92.73376, 91.27863, 89.15242, 89.31269, 
    91.05988, 92.17466, 91.37316, 91.41622, 92.72636, 94.31723,
  92.37487, 92.17799, 91.41553, 90.4892, 90.00282, 89.10106, 87.04726, 
    84.81566, 82.27917, 79.78806, 74.15566, 68.09465, 64.61887, 64.36955, 
    66.42295, 69.61932, 73.69915, 80.02668, 86.2827, 88.02354,
  80.78298, 80.45201, 79.41755, 77.19287, 74.21328, 70.90347, 68.3314, 
    67.25011, 66.53024, 66.63924, 65.926, 65.46037, 66.2202, 68.19367, 
    70.01898, 70.74322, 70.28625, 70.23486, 70.74574, 70.54175,
  79.27809, 79.03497, 77.76959, 75.15334, 71.25109, 68.02479, 65.255, 
    63.87289, 63.64126, 64.60026, 65.54762, 67.19524, 69.5436, 71.86909, 
    73.01209, 73.62477, 73.43317, 73.13465, 73.30375, 74.42599,
  76.81366, 77.47233, 75.62317, 71.47828, 66.47199, 63.4263, 61.94608, 
    61.67241, 62.23563, 63.82353, 66.72684, 70.37658, 73.5173, 75.48281, 
    75.76226, 75.74701, 74.84489, 73.66897, 73.68858, 74.68499,
  71.05982, 69.08096, 65.1989, 60.95345, 57.91884, 57.03664, 57.73422, 
    58.82198, 60.35466, 62.76599, 66.06871, 69.69015, 72.69817, 74.61146, 
    75.07155, 74.67497, 72.52214, 70.13746, 68.13469, 66.70573,
  62.19204, 57.83405, 55.80669, 55.62794, 56.30608, 57.73314, 58.83397, 
    58.23901, 57.00458, 57.17825, 58.94392, 61.49005, 64.32321, 66.93961, 
    69.4767, 70.19569, 67.43777, 63.70792, 61.43116, 60.55825,
  60.00661, 60.75495, 62.08223, 64.46676, 66.27565, 65.65942, 62.55649, 
    60.7638, 59.57166, 56.9856, 56.38796, 58.04719, 60.64682, 62.69976, 
    64.55711, 65.05193, 63.93134, 62.36448, 61.59513, 62.16031,
  66.79579, 68.18753, 69.41352, 70.35666, 68.83643, 66.82329, 66.16498, 
    68.64828, 69.73102, 65.72814, 60.79543, 60.89844, 66.94974, 68.74442, 
    68.26937, 67.64861, 67.0584, 66.31132, 65.99249, 66.99352,
  88.609, 88.9129, 89.35703, 89.58056, 89.88323, 90.31568, 90.47955, 
    90.59157, 89.16118, 89.41843, 89.58453, 89.66906, 89.76942, 89.92445, 
    90.09928, 90.19556, 89.3242, 89.37884, 89.41559, 89.4796,
  83.50027, 84.45282, 85.40108, 86.38496, 87.47705, 88.68792, 89.89538, 
    91.12411, 87.74897, 88.90193, 89.69777, 90.41906, 90.98679, 91.55551, 
    92.28655, 93.00558, 91.22588, 91.55207, 91.84856, 92.22795,
  85.09618, 86.47843, 87.49725, 88.23017, 89.37714, 90.60735, 91.88024, 
    93.13723, 89.11244, 90.08474, 90.72935, 91.42802, 91.84574, 92.1894, 
    92.48628, 92.92882, 91.36217, 91.64245, 91.75526, 91.90024,
  85.69303, 87.26197, 88.94791, 90.5173, 91.41416, 92.21964, 92.95592, 
    93.63611, 90.9937, 91.25299, 91.27473, 92.05956, 93.35052, 94.11979, 
    94.81309, 95.22103, 95.74983, 95.27264, 94.45729, 93.45393,
  84.85725, 86.04678, 86.42396, 85.67586, 86.85174, 87.73362, 88.45018, 
    88.91193, 87.94398, 88.42483, 89.46203, 90.39451, 91.30072, 92.28681, 
    93.16993, 93.60343, 96.98302, 96.74683, 96.36903, 95.66586,
  82.56306, 83.56171, 84.13232, 84.87933, 85.47791, 85.95991, 86.00638, 
    85.72562, 80.97152, 81.09812, 81.47396, 82.24639, 83.32902, 84.48576, 
    85.66669, 86.7346, 94.13512, 94.68295, 94.95634, 94.61739,
  93.54938, 90.57149, 87.96381, 87.17788, 87.76167, 87.61079, 87.19888, 
    86.53236, 79.53448, 80.37038, 80.28065, 74.30634, 76.56163, 83.89491, 
    85.50579, 81.93359, 89.03914, 91.28963, 93.061, 93.67842,
  97.15588, 96.2106, 94.53758, 93.2066, 93.91686, 93.86451, 93.88658, 
    93.46226, 89.66816, 89.51099, 87.47245, 88.26347, 89.96706, 93.91555, 
    94.9223, 85.15292, 94.1926, 93.46297, 91.64505, 92.47969,
  96.58619, 96.36151, 95.48752, 94.63628, 93.82732, 93.34805, 93.19348, 
    93.28653, 92.12846, 93.00917, 93.56448, 93.34886, 93.48616, 93.77395, 
    94.44027, 95.70678, 95.87537, 97.45126, 96.9576, 97.33305,
  95.90493, 95.88762, 95.74536, 95.89227, 95.49886, 94.83835, 94.71727, 
    94.84889, 94.38562, 94.72091, 94.90517, 94.92635, 93.89286, 92.894, 
    93.7248, 94.85355, 95.51345, 96.22449, 96.81009, 97.11147,
  95.80334, 95.73128, 95.72832, 95.75616, 95.35781, 94.94672, 95.06435, 
    95.32649, 95.15401, 95.09362, 94.99785, 94.84078, 94.25739, 93.93702, 
    93.40908, 93.45232, 93.33428, 93.61575, 94.03213, 94.36234,
  95.87843, 95.70851, 95.27673, 94.78841, 94.27863, 94.36084, 94.58128, 
    94.77731, 94.40265, 94.5924, 93.84163, 92.76368, 92.33602, 92.48273, 
    91.98473, 91.85608, 91.22127, 91.49603, 92.55194, 93.16766,
  94.16338, 94.41628, 94.5695, 94.33678, 94.04425, 93.39246, 92.17838, 
    90.91929, 89.97933, 89.00486, 85.57747, 78.02666, 74.21856, 73.92089, 
    74.40086, 76.01141, 79.06516, 82.58479, 85.38322, 86.80526,
  86.74515, 86.96786, 87.3227, 85.90944, 81.47916, 76.54398, 72.23557, 
    70.03638, 68.89806, 68.8157, 67.59385, 66.31068, 66.57243, 68.44991, 
    70.90773, 72.71643, 73.9437, 75.30574, 77.17347, 79.30849,
  84.4836, 84.19073, 82.49574, 79.36344, 74.76008, 71.54102, 69.25411, 
    67.83772, 67.73102, 69.04715, 70.28819, 71.63869, 73.54847, 75.61906, 
    77.08699, 77.4763, 77.15446, 77.15075, 78.26665, 81.11185,
  80.74612, 81.14505, 78.70613, 73.83881, 68.98478, 66.69609, 66.17759, 
    66.70178, 67.90977, 70.00713, 72.47179, 75.57169, 78.54701, 80.76289, 
    80.6255, 79.91996, 79.42898, 78.60263, 79.13939, 81.18186,
  76.20496, 74.24358, 70.39124, 65.85323, 63.64817, 63.03072, 62.95248, 
    63.97334, 65.41827, 67.85667, 70.5882, 74.01851, 77.63241, 80.05271, 
    80.06287, 79.35762, 78.11939, 76.79914, 76.42435, 76.87436,
  69.15688, 66.03324, 64.74166, 63.46961, 62.55168, 62.05645, 61.84727, 
    60.9156, 59.02358, 58.81698, 59.75974, 62.39579, 66.51761, 69.93262, 
    72.04633, 72.73006, 71.04943, 68.67365, 67.81168, 69.082,
  65.18978, 66.71393, 68.28641, 68.85825, 67.65556, 64.9138, 60.98755, 
    57.90487, 54.43315, 51.18723, 50.59245, 52.65274, 55.98347, 58.56968, 
    60.9522, 62.2267, 62.80406, 62.926, 63.94051, 66.85204,
  68.17101, 69.26753, 70.16818, 69.73458, 67.22097, 63.44703, 60.49933, 
    59.94702, 58.25105, 53.96359, 50.21961, 51.82551, 58.37508, 61.8357, 
    62.88547, 63.70344, 65.37298, 67.26636, 69.90611, 73.22445,
  89.12636, 89.4614, 89.73013, 90.08813, 90.49535, 90.90154, 91.30602, 
    91.63762, 90.16696, 90.46536, 90.77396, 91.06967, 91.31654, 91.60416, 
    91.82911, 92.16157, 91.41087, 91.58636, 91.75822, 92.0507,
  85.69506, 86.4969, 87.31724, 88.21929, 89.1537, 90.02069, 90.91573, 
    91.85177, 88.34193, 89.21027, 89.99326, 90.75661, 91.48685, 92.22185, 
    92.99342, 93.79789, 92.04114, 92.71863, 93.2965, 93.90443,
  85.0059, 85.9136, 87.03998, 88.28199, 89.42886, 90.75167, 91.9587, 
    93.46645, 89.41599, 90.62556, 91.50703, 92.31778, 93.22275, 94.17249, 
    95.13268, 95.97668, 94.30376, 94.84152, 95.25953, 95.32898,
  85.60783, 87.1151, 88.73589, 90.31673, 91.90896, 93.37848, 94.7055, 
    95.70452, 93.33681, 94.11471, 94.64704, 94.95362, 95.11736, 95.18666, 
    95.61439, 95.71722, 96.51637, 96.38905, 96.48267, 96.13758,
  84.89723, 87.2158, 89.17696, 90.73365, 92.32804, 93.52126, 94.43604, 
    95.14668, 94.05721, 94.4491, 94.24294, 94.0315, 94.18307, 94.3947, 
    94.601, 94.56442, 98.27877, 98.22531, 98.0214, 97.58329,
  85.35185, 87.57565, 89.59953, 91.25391, 92.45763, 93.15097, 93.70103, 
    93.95906, 89.39124, 89.27857, 89.2146, 89.64468, 90.27628, 91.23914, 
    92.39287, 93.45592, 98.77247, 98.9912, 98.9409, 98.60909,
  90.96671, 88.95423, 88.33873, 89.1646, 89.85364, 89.4952, 89.20425, 
    89.07461, 81.72141, 81.3737, 79.73669, 78.98242, 81.09166, 87.54227, 
    87.02039, 87.64054, 95.34365, 97.37656, 98.32056, 98.55834,
  92.12396, 91.71731, 91.66611, 91.82751, 92.13261, 91.57689, 91.58893, 
    91.29268, 86.8933, 85.071, 80.35474, 85.14971, 87.37561, 92.70294, 
    89.11998, 84.07039, 89.66982, 94.57336, 94.15179, 96.17076,
  93.67297, 93.10026, 91.91206, 91.17325, 90.94757, 90.69505, 90.55582, 
    90.46128, 88.38421, 88.19518, 87.97022, 88.04433, 89.64313, 91.34264, 
    93.09979, 94.25278, 94.34208, 95.28682, 94.71233, 95.80148,
  95.36063, 95.46169, 95.55, 94.86865, 94.65484, 94.58582, 94.24242, 
    94.08227, 93.95758, 93.76926, 93.46625, 93.1393, 93.34606, 93.8012, 
    94.31777, 95.63311, 96.41074, 96.72069, 96.62096, 96.32957,
  95.48937, 95.47292, 95.57552, 95.8564, 95.84338, 95.85989, 95.5125, 
    95.41924, 95.54803, 95.57485, 95.03793, 94.75723, 94.33324, 94.22587, 
    94.26043, 95.03274, 95.60491, 95.19999, 94.87977, 94.58964,
  94.33001, 94.45174, 94.35564, 94.19715, 94.39539, 94.26285, 94.09069, 
    94.30093, 94.40318, 94.41055, 94.16878, 93.77896, 93.24632, 93.024, 
    93.51138, 93.97529, 94.33997, 94.46935, 94.39352, 94.33096,
  88.64445, 89.12266, 89.48273, 89.98489, 90.66469, 90.18948, 88.6783, 
    87.90173, 88.14387, 88.0686, 87.14576, 85.59967, 84.68818, 85.51276, 
    87.20138, 88.15849, 87.93333, 87.83617, 88.23782, 89.27096,
  84.90213, 85.43855, 86.00737, 85.43637, 82.83469, 79.2315, 75.97392, 
    74.22888, 74.33865, 75.82793, 76.50627, 76.52354, 77.00267, 78.71989, 
    81.05069, 81.77783, 81.29063, 82.08588, 83.82008, 85.73005,
  85.40762, 86.51618, 86.96132, 85.37651, 81.22579, 77.46445, 74.64709, 
    73.1145, 73.16389, 75.06313, 77.49453, 79.88705, 81.67218, 83.15096, 
    84.08208, 84.03651, 82.94983, 82.38705, 83.12579, 85.3443,
  83.21449, 84.42175, 83.65591, 80.31356, 76.08496, 74.14221, 73.88336, 
    74.23907, 75.98573, 78.70048, 81.61548, 83.98601, 85.53611, 86.62379, 
    86.16817, 84.92745, 83.13875, 81.40516, 81.17575, 82.07327,
  80.11454, 79.27293, 76.59651, 73.4086, 71.93156, 73.21077, 74.72791, 
    75.76893, 77.26123, 78.91931, 80.45676, 82.34642, 84.14986, 85.09487, 
    84.34818, 82.30523, 79.29346, 76.50311, 74.52405, 73.79091,
  74.46515, 71.88083, 70.97222, 71.93839, 73.25758, 74.67936, 75.4819, 
    74.0758, 70.7289, 69.52139, 70.20005, 72.26597, 74.66635, 75.94512, 
    76.4346, 75.64117, 72.51921, 69.00674, 67.16875, 67.38728,
  71.39501, 73.29038, 75.00249, 75.76629, 75.89171, 74.44814, 71.42114, 
    67.09987, 62.67251, 59.48172, 58.93935, 60.68055, 63.95771, 67.14864, 
    68.93729, 69.06831, 68.39293, 67.58773, 67.59353, 68.30827,
  72.32693, 73.78093, 73.10394, 72.04498, 71.23317, 69.56831, 67.23677, 
    63.43821, 63.92851, 62.26643, 60.17223, 61.05844, 67.29062, 71.2075, 
    70.97546, 70.17451, 69.70806, 70.31026, 71.31174, 71.96861,
  91.44809, 91.66164, 91.81742, 91.98062, 92.01276, 92.00135, 92.13506, 
    92.19342, 90.77084, 90.76516, 90.96467, 91.05332, 91.1897, 91.32604, 
    91.40299, 91.48151, 90.54983, 90.57541, 90.60886, 90.69357,
  85.24937, 85.48785, 85.99204, 86.43094, 86.9384, 87.58467, 88.57504, 
    89.11788, 86.17255, 87.03139, 87.7996, 88.37601, 89.0016, 89.63566, 
    90.05051, 90.46011, 88.35456, 88.60172, 88.9237, 89.3385,
  81.12431, 81.79145, 82.62906, 83.18066, 84.18713, 85.35401, 86.44003, 
    87.64559, 83.91792, 85.10661, 86.24564, 87.54995, 88.78102, 89.70271, 
    90.27992, 91.1144, 89.29219, 89.5969, 89.95528, 90.23089,
  80.9297, 81.60825, 82.33701, 83.26079, 84.05903, 85.23982, 86.37723, 
    87.47364, 85.01184, 85.74561, 86.68483, 87.52085, 88.57964, 88.96327, 
    89.15256, 89.25525, 89.92667, 89.41711, 89.56737, 89.43054,
  80.43243, 82.82311, 84.75478, 86.36188, 88.08858, 89.19492, 90.13615, 
    90.92628, 89.67474, 89.88817, 89.92721, 90.32404, 90.22188, 90.33604, 
    90.34371, 90.25446, 94.90108, 94.37499, 93.40989, 92.55029,
  79.87, 82.67743, 85.02766, 86.26923, 87.29717, 88.29794, 88.90195, 
    89.00178, 85.1427, 85.46175, 85.97768, 86.80894, 87.46559, 88.52172, 
    89.81921, 91.12234, 97.60638, 97.78215, 97.73178, 97.39719,
  87.93222, 83.60091, 82.85329, 84.01416, 84.41905, 84.23631, 83.99754, 
    83.80155, 75.77188, 74.47368, 72.97333, 74.98318, 76.69712, 81.3893, 
    82.19207, 85.57985, 93.35909, 95.63696, 96.80153, 97.29794,
  89.75894, 90.26264, 91.42225, 92.5764, 92.67274, 92.11102, 91.42975, 
    90.82169, 82.88423, 79.09122, 74.91882, 80.31293, 82.14307, 88.54573, 
    80.22871, 77.76046, 79.15327, 91.58929, 90.69492, 92.74844,
  90.62286, 90.09777, 90.41944, 91.4126, 91.83208, 91.92006, 91.56749, 
    90.91813, 87.62701, 86.92293, 86.47465, 85.94659, 85.62832, 85.43887, 
    87.19572, 90.19321, 91.97924, 91.60905, 92.5863, 94.78312,
  93.38673, 93.16024, 93.28277, 94.21758, 94.66365, 94.47284, 94.42598, 
    94.17593, 92.54395, 90.83896, 90.66453, 90.31806, 89.82665, 89.05578, 
    88.30283, 89.30795, 91.33284, 93.52869, 94.97649, 95.61607,
  91.07861, 91.35603, 91.3896, 91.72186, 92.11106, 92.68369, 93.38113, 
    93.64973, 93.73654, 93.67008, 93.90296, 94.18099, 93.96429, 92.81234, 
    90.21255, 88.14841, 86.85229, 86.90884, 88.59177, 90.27828,
  87.82471, 88.01861, 88.25435, 88.78571, 89.3428, 89.59425, 89.59976, 
    89.65371, 89.37206, 88.54897, 88.61231, 90.08528, 92.00015, 93.30373, 
    93.70888, 92.61208, 90.07843, 88.09201, 87.20648, 87.71262,
  85.86485, 85.95393, 86.33294, 86.82038, 87.33516, 86.78876, 85.96225, 
    85.52868, 84.8943, 83.83492, 82.4426, 82.40176, 84.30611, 87.1742, 
    88.98733, 90.04581, 89.93927, 89.39529, 88.90865, 88.87407,
  87.11257, 86.95045, 87.13309, 86.61064, 84.85566, 82.42012, 80.78365, 
    80.29518, 80.76437, 81.82693, 81.45129, 80.60843, 80.08038, 81.4576, 
    83.89008, 85.37902, 85.08916, 86.01255, 87.49905, 88.82468,
  87.86531, 87.98333, 87.86685, 86.08907, 82.51519, 80.26978, 79.41601, 
    79.2778, 79.92186, 81.49277, 83.09648, 84.216, 83.98283, 83.39529, 
    83.74914, 84.23751, 83.67759, 83.71537, 84.93969, 87.4865,
  86.00185, 86.50753, 84.91483, 81.32465, 77.867, 76.77679, 77.5079, 
    78.76208, 80.04148, 82.12397, 84.59582, 86.46084, 86.94716, 86.49524, 
    85.67841, 84.98366, 83.6435, 82.8194, 83.62476, 84.85889,
  83.51066, 82.53691, 80.0031, 77.42001, 76.20304, 77.06575, 78.9127, 
    79.99328, 80.38633, 81.67112, 83.48209, 84.82047, 85.35446, 85.32668, 
    84.60071, 83.68895, 81.70484, 79.60397, 78.11585, 76.9676,
  80.27482, 78.06759, 77.14984, 78.04604, 79.50267, 80.69393, 81.08243, 
    79.14809, 73.99506, 71.88085, 72.83691, 75.27429, 77.5179, 78.91724, 
    79.20642, 78.70898, 76.1686, 72.92442, 70.57545, 69.61903,
  78.69959, 79.60489, 81.61304, 82.84615, 83.28924, 81.59545, 77.40047, 
    69.99107, 62.72016, 59.24093, 59.89368, 63.16311, 67.00726, 69.86009, 
    71.28391, 71.82669, 70.98501, 70.24709, 70.12183, 70.55403,
  78.56296, 79.19095, 78.90386, 78.00187, 76.5765, 73.66414, 69.25168, 
    63.40796, 63.06129, 63.01234, 64.50167, 66.44123, 71.52995, 74.49757, 
    74.53848, 74.47372, 73.41979, 73.30776, 73.84573, 74.36893 ;
}
