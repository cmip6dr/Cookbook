netcdf zsatcalc_Omon_exAA07_abrupt4xCO2_r1i1p1_013601-014012_box {
dimensions:
	x = 20 ;
	y = 20 ;
	nv4 = 4 ;
	time = UNLIMITED ; // (4 currently)
	bnds = 2 ;
variables:
	float lon(y, x) ;
		lon:standard_name = "longitude" ;
		lon:long_name = "longitude coordinate" ;
		lon:units = "degrees_east" ;
		lon:_CoordinateAxisType = "Lon" ;
		lon:bounds = "lon_bnds" ;
	float lon_bnds(y, x, nv4) ;
	float lat(y, x) ;
		lat:standard_name = "latitude" ;
		lat:long_name = "latitude coordinate" ;
		lat:units = "degrees_north" ;
		lat:_CoordinateAxisType = "Lat" ;
		lat:bounds = "lat_bnds" ;
	float lat_bnds(y, x, nv4) ;
	double time(time) ;
		time:standard_name = "time" ;
		time:long_name = "time" ;
		time:bounds = "time_bnds" ;
		time:units = "days since 1-1-1 00:00:00" ;
		time:calendar = "365_day" ;
		time:axis = "T" ;
	double time_bnds(time, bnds) ;
	double average_DT(time) ;
		average_DT:long_name = "Length of average period" ;
		average_DT:units = "days" ;
	float zsatcalc(time, y, x) ;
		zsatcalc:standard_name = "minimum_depth_of_calcite_undersaturation_in_sea_water" ;
		zsatcalc:long_name = "Calcite Saturation Depth" ;
		zsatcalc:units = "m" ;
		zsatcalc:coordinates = "lat lon" ;
		zsatcalc:_FillValue = 1.e+20f ;
		zsatcalc:missing_value = 1.e+20f ;
		zsatcalc:cell_methods = "time: mean area: where sea" ;
		zsatcalc:comments = "Note: This model output is presented on the model\'s tripolar grid. The North Pole singularity is avoided by using this nonregular grid north of 65N. More information about the ocean and sea ice model\'s grid can be found at http://nomads.gfdl.noaa.gov/." ;
		zsatcalc:original_name = "zsatcalc" ;
		zsatcalc:original_units = "m" ;
		zsatcalc:associated_files = "baseURL: http://cmip-pcmdi.llnl.gov/CMIP5/dataLocation gridspecFile: gridspec_ocnBgchem_fx_GFDL-ESM2M_abrupt4xCO2_r0i0p0.nc areacello: areacello_fx_GFDL-ESM2M_abrupt4xCO2_r0i0p0.nc" ;

// global attributes:
		:CDI = "Climate Data Interface version ?? (http://mpimet.mpg.de/cdi)" ;
		:Conventions = "CF-1.4" ;
		:history = "reset by cdo to create anonymous sample file" ;
		:source = "201707_compliance_checker_evaluation/work/p1.py" ;
		:institution = "CEDA" ;
		:title = "Dummy file with known metadata errors" ;
		:institute_id = "CEDA" ;
		:contact = "none" ;
		:project_id = "CMIP5" ;
		:table_id = "Table Omon (31 Jan 2011)" ;
		:experiment_id = "abrupt4xCO2" ;
		:realization = 1 ;
		:modeling_realm = "ocnBgchem" ;
		:tracking_id = "431d6e16-bd03-42ed-ad62-15c7f90621e8" ;
		:references = "The GFDL Data Portal (http://nomads.gfdl.noaa.gov/) provides access to NOAA/GFDL\'s publicly available model input and output data sets. From this web site one can view and download data sets and documentation, including those related to the GFDL coupled models experiments run for the IPCC\'s 5th Assessment Report and the US CCSP." ;
		:comment = "this is a sample file with known metadata errors" ;
		:gfdl_experiment_name = "ESM2M-C1_abrupt-4xco2_S1" ;
		:creation_date = "2012-02-02T17:54:27Z" ;
		:model_id = "exAA07" ;
		:branch_time = "0.0" ;
		:experiment = "abrupt 4XCO2" ;
		:forcing = "GHG (GHG includes only time varying CO2)" ;
		:frequency = "mon" ;
		:initialization_method = 1 ;
		:parent_experiment_id = "N/A" ;
		:physics_version = 1 ;
		:product = "output1" ;
		:parent_experiment_rip = "N/A" ;
		:CDO = "Climate Data Operators version 1.7.0 (http://mpimet.mpg.de/cdo)" ;
data:

 lon =
  -279.5, -278.5, -277.5, -276.5, -275.5, -274.5, -273.5, -272.5, -271.5, 
    -270.5, -269.5, -268.5, -267.5, -266.5, -265.5, -264.5, -263.5, -262.5, 
    -261.5, -260.5,
  -279.5, -278.5, -277.5, -276.5, -275.5, -274.5, -273.5, -272.5, -271.5, 
    -270.5, -269.5, -268.5, -267.5, -266.5, -265.5, -264.5, -263.5, -262.5, 
    -261.5, -260.5,
  -279.5, -278.5, -277.5, -276.5, -275.5, -274.5, -273.5, -272.5, -271.5, 
    -270.5, -269.5, -268.5, -267.5, -266.5, -265.5, -264.5, -263.5, -262.5, 
    -261.5, -260.5,
  -279.5, -278.5, -277.5, -276.5, -275.5, -274.5, -273.5, -272.5, -271.5, 
    -270.5, -269.5, -268.5, -267.5, -266.5, -265.5, -264.5, -263.5, -262.5, 
    -261.5, -260.5,
  -279.5, -278.5, -277.5, -276.5, -275.5, -274.5, -273.5, -272.5, -271.5, 
    -270.5, -269.5, -268.5, -267.5, -266.5, -265.5, -264.5, -263.5, -262.5, 
    -261.5, -260.5,
  -279.5, -278.5, -277.5, -276.5, -275.5, -274.5, -273.5, -272.5, -271.5, 
    -270.5, -269.5, -268.5, -267.5, -266.5, -265.5, -264.5, -263.5, -262.5, 
    -261.5, -260.5,
  -279.5, -278.5, -277.5, -276.5, -275.5, -274.5, -273.5, -272.5, -271.5, 
    -270.5, -269.5, -268.5, -267.5, -266.5, -265.5, -264.5, -263.5, -262.5, 
    -261.5, -260.5,
  -279.5, -278.5, -277.5, -276.5, -275.5, -274.5, -273.5, -272.5, -271.5, 
    -270.5, -269.5, -268.5, -267.5, -266.5, -265.5, -264.5, -263.5, -262.5, 
    -261.5, -260.5,
  -279.5, -278.5, -277.5, -276.5, -275.5, -274.5, -273.5, -272.5, -271.5, 
    -270.5, -269.5, -268.5, -267.5, -266.5, -265.5, -264.5, -263.5, -262.5, 
    -261.5, -260.5,
  -279.5, -278.5, -277.5, -276.5, -275.5, -274.5, -273.5, -272.5, -271.5, 
    -270.5, -269.5, -268.5, -267.5, -266.5, -265.5, -264.5, -263.5, -262.5, 
    -261.5, -260.5,
  -279.5, -278.5, -277.5, -276.5, -275.5, -274.5, -273.5, -272.5, -271.5, 
    -270.5, -269.5, -268.5, -267.5, -266.5, -265.5, -264.5, -263.5, -262.5, 
    -261.5, -260.5,
  -279.5, -278.5, -277.5, -276.5, -275.5, -274.5, -273.5, -272.5, -271.5, 
    -270.5, -269.5, -268.5, -267.5, -266.5, -265.5, -264.5, -263.5, -262.5, 
    -261.5, -260.5,
  -279.5, -278.5, -277.5, -276.5, -275.5, -274.5, -273.5, -272.5, -271.5, 
    -270.5, -269.5, -268.5, -267.5, -266.5, -265.5, -264.5, -263.5, -262.5, 
    -261.5, -260.5,
  -279.5, -278.5, -277.5, -276.5, -275.5, -274.5, -273.5, -272.5, -271.5, 
    -270.5, -269.5, -268.5, -267.5, -266.5, -265.5, -264.5, -263.5, -262.5, 
    -261.5, -260.5,
  -279.5, -278.5, -277.5, -276.5, -275.5, -274.5, -273.5, -272.5, -271.5, 
    -270.5, -269.5, -268.5, -267.5, -266.5, -265.5, -264.5, -263.5, -262.5, 
    -261.5, -260.5,
  -279.5, -278.5, -277.5, -276.5, -275.5, -274.5, -273.5, -272.5, -271.5, 
    -270.5, -269.5, -268.5, -267.5, -266.5, -265.5, -264.5, -263.5, -262.5, 
    -261.5, -260.5,
  -279.5, -278.5, -277.5, -276.5, -275.5, -274.5, -273.5, -272.5, -271.5, 
    -270.5, -269.5, -268.5, -267.5, -266.5, -265.5, -264.5, -263.5, -262.5, 
    -261.5, -260.5,
  -279.5, -278.5, -277.5, -276.5, -275.5, -274.5, -273.5, -272.5, -271.5, 
    -270.5, -269.5, -268.5, -267.5, -266.5, -265.5, -264.5, -263.5, -262.5, 
    -261.5, -260.5,
  -279.5, -278.5, -277.5, -276.5, -275.5, -274.5, -273.5, -272.5, -271.5, 
    -270.5, -269.5, -268.5, -267.5, -266.5, -265.5, -264.5, -263.5, -262.5, 
    -261.5, -260.5,
  -279.5, -278.5, -277.5, -276.5, -275.5, -274.5, -273.5, -272.5, -271.5, 
    -270.5, -269.5, -268.5, -267.5, -266.5, -265.5, -264.5, -263.5, -262.5, 
    -261.5, -260.5 ;

 lon_bnds =
  -280, -279, -279, -280,
  -279, -278, -278, -279,
  -278, -277, -277, -278,
  -277, -276, -276, -277,
  -276, -275, -275, -276,
  -275, -274, -274, -275,
  -274, -273, -273, -274,
  -273, -272, -272, -273,
  -272, -271, -271, -272,
  -271, -270, -270, -271,
  -270, -269, -269, -270,
  -269, -268, -268, -269,
  -268, -267, -267, -268,
  -267, -266, -266, -267,
  -266, -265, -265, -266,
  -265, -264, -264, -265,
  -264, -263, -263, -264,
  -263, -262, -262, -263,
  -262, -261, -261, -262,
  -261, -260, -260, -261,
  -280, -279, -279, -280,
  -279, -278, -278, -279,
  -278, -277, -277, -278,
  -277, -276, -276, -277,
  -276, -275, -275, -276,
  -275, -274, -274, -275,
  -274, -273, -273, -274,
  -273, -272, -272, -273,
  -272, -271, -271, -272,
  -271, -270, -270, -271,
  -270, -269, -269, -270,
  -269, -268, -268, -269,
  -268, -267, -267, -268,
  -267, -266, -266, -267,
  -266, -265, -265, -266,
  -265, -264, -264, -265,
  -264, -263, -263, -264,
  -263, -262, -262, -263,
  -262, -261, -261, -262,
  -261, -260, -260, -261,
  -280, -279, -279, -280,
  -279, -278, -278, -279,
  -278, -277, -277, -278,
  -277, -276, -276, -277,
  -276, -275, -275, -276,
  -275, -274, -274, -275,
  -274, -273, -273, -274,
  -273, -272, -272, -273,
  -272, -271, -271, -272,
  -271, -270, -270, -271,
  -270, -269, -269, -270,
  -269, -268, -268, -269,
  -268, -267, -267, -268,
  -267, -266, -266, -267,
  -266, -265, -265, -266,
  -265, -264, -264, -265,
  -264, -263, -263, -264,
  -263, -262, -262, -263,
  -262, -261, -261, -262,
  -261, -260, -260, -261,
  -280, -279, -279, -280,
  -279, -278, -278, -279,
  -278, -277, -277, -278,
  -277, -276, -276, -277,
  -276, -275, -275, -276,
  -275, -274, -274, -275,
  -274, -273, -273, -274,
  -273, -272, -272, -273,
  -272, -271, -271, -272,
  -271, -270, -270, -271,
  -270, -269, -269, -270,
  -269, -268, -268, -269,
  -268, -267, -267, -268,
  -267, -266, -266, -267,
  -266, -265, -265, -266,
  -265, -264, -264, -265,
  -264, -263, -263, -264,
  -263, -262, -262, -263,
  -262, -261, -261, -262,
  -261, -260, -260, -261,
  -280, -279, -279, -280,
  -279, -278, -278, -279,
  -278, -277, -277, -278,
  -277, -276, -276, -277,
  -276, -275, -275, -276,
  -275, -274, -274, -275,
  -274, -273, -273, -274,
  -273, -272, -272, -273,
  -272, -271, -271, -272,
  -271, -270, -270, -271,
  -270, -269, -269, -270,
  -269, -268, -268, -269,
  -268, -267, -267, -268,
  -267, -266, -266, -267,
  -266, -265, -265, -266,
  -265, -264, -264, -265,
  -264, -263, -263, -264,
  -263, -262, -262, -263,
  -262, -261, -261, -262,
  -261, -260, -260, -261,
  -280, -279, -279, -280,
  -279, -278, -278, -279,
  -278, -277, -277, -278,
  -277, -276, -276, -277,
  -276, -275, -275, -276,
  -275, -274, -274, -275,
  -274, -273, -273, -274,
  -273, -272, -272, -273,
  -272, -271, -271, -272,
  -271, -270, -270, -271,
  -270, -269, -269, -270,
  -269, -268, -268, -269,
  -268, -267, -267, -268,
  -267, -266, -266, -267,
  -266, -265, -265, -266,
  -265, -264, -264, -265,
  -264, -263, -263, -264,
  -263, -262, -262, -263,
  -262, -261, -261, -262,
  -261, -260, -260, -261,
  -280, -279, -279, -280,
  -279, -278, -278, -279,
  -278, -277, -277, -278,
  -277, -276, -276, -277,
  -276, -275, -275, -276,
  -275, -274, -274, -275,
  -274, -273, -273, -274,
  -273, -272, -272, -273,
  -272, -271, -271, -272,
  -271, -270, -270, -271,
  -270, -269, -269, -270,
  -269, -268, -268, -269,
  -268, -267, -267, -268,
  -267, -266, -266, -267,
  -266, -265, -265, -266,
  -265, -264, -264, -265,
  -264, -263, -263, -264,
  -263, -262, -262, -263,
  -262, -261, -261, -262,
  -261, -260, -260, -261,
  -280, -279, -279, -280,
  -279, -278, -278, -279,
  -278, -277, -277, -278,
  -277, -276, -276, -277,
  -276, -275, -275, -276,
  -275, -274, -274, -275,
  -274, -273, -273, -274,
  -273, -272, -272, -273,
  -272, -271, -271, -272,
  -271, -270, -270, -271,
  -270, -269, -269, -270,
  -269, -268, -268, -269,
  -268, -267, -267, -268,
  -267, -266, -266, -267,
  -266, -265, -265, -266,
  -265, -264, -264, -265,
  -264, -263, -263, -264,
  -263, -262, -262, -263,
  -262, -261, -261, -262,
  -261, -260, -260, -261,
  -280, -279, -279, -280,
  -279, -278, -278, -279,
  -278, -277, -277, -278,
  -277, -276, -276, -277,
  -276, -275, -275, -276,
  -275, -274, -274, -275,
  -274, -273, -273, -274,
  -273, -272, -272, -273,
  -272, -271, -271, -272,
  -271, -270, -270, -271,
  -270, -269, -269, -270,
  -269, -268, -268, -269,
  -268, -267, -267, -268,
  -267, -266, -266, -267,
  -266, -265, -265, -266,
  -265, -264, -264, -265,
  -264, -263, -263, -264,
  -263, -262, -262, -263,
  -262, -261, -261, -262,
  -261, -260, -260, -261,
  -280, -279, -279, -280,
  -279, -278, -278, -279,
  -278, -277, -277, -278,
  -277, -276, -276, -277,
  -276, -275, -275, -276,
  -275, -274, -274, -275,
  -274, -273, -273, -274,
  -273, -272, -272, -273,
  -272, -271, -271, -272,
  -271, -270, -270, -271,
  -270, -269, -269, -270,
  -269, -268, -268, -269,
  -268, -267, -267, -268,
  -267, -266, -266, -267,
  -266, -265, -265, -266,
  -265, -264, -264, -265,
  -264, -263, -263, -264,
  -263, -262, -262, -263,
  -262, -261, -261, -262,
  -261, -260, -260, -261,
  -280, -279, -279, -280,
  -279, -278, -278, -279,
  -278, -277, -277, -278,
  -277, -276, -276, -277,
  -276, -275, -275, -276,
  -275, -274, -274, -275,
  -274, -273, -273, -274,
  -273, -272, -272, -273,
  -272, -271, -271, -272,
  -271, -270, -270, -271,
  -270, -269, -269, -270,
  -269, -268, -268, -269,
  -268, -267, -267, -268,
  -267, -266, -266, -267,
  -266, -265, -265, -266,
  -265, -264, -264, -265,
  -264, -263, -263, -264,
  -263, -262, -262, -263,
  -262, -261, -261, -262,
  -261, -260, -260, -261,
  -280, -279, -279, -280,
  -279, -278, -278, -279,
  -278, -277, -277, -278,
  -277, -276, -276, -277,
  -276, -275, -275, -276,
  -275, -274, -274, -275,
  -274, -273, -273, -274,
  -273, -272, -272, -273,
  -272, -271, -271, -272,
  -271, -270, -270, -271,
  -270, -269, -269, -270,
  -269, -268, -268, -269,
  -268, -267, -267, -268,
  -267, -266, -266, -267,
  -266, -265, -265, -266,
  -265, -264, -264, -265,
  -264, -263, -263, -264,
  -263, -262, -262, -263,
  -262, -261, -261, -262,
  -261, -260, -260, -261,
  -280, -279, -279, -280,
  -279, -278, -278, -279,
  -278, -277, -277, -278,
  -277, -276, -276, -277,
  -276, -275, -275, -276,
  -275, -274, -274, -275,
  -274, -273, -273, -274,
  -273, -272, -272, -273,
  -272, -271, -271, -272,
  -271, -270, -270, -271,
  -270, -269, -269, -270,
  -269, -268, -268, -269,
  -268, -267, -267, -268,
  -267, -266, -266, -267,
  -266, -265, -265, -266,
  -265, -264, -264, -265,
  -264, -263, -263, -264,
  -263, -262, -262, -263,
  -262, -261, -261, -262,
  -261, -260, -260, -261,
  -280, -279, -279, -280,
  -279, -278, -278, -279,
  -278, -277, -277, -278,
  -277, -276, -276, -277,
  -276, -275, -275, -276,
  -275, -274, -274, -275,
  -274, -273, -273, -274,
  -273, -272, -272, -273,
  -272, -271, -271, -272,
  -271, -270, -270, -271,
  -270, -269, -269, -270,
  -269, -268, -268, -269,
  -268, -267, -267, -268,
  -267, -266, -266, -267,
  -266, -265, -265, -266,
  -265, -264, -264, -265,
  -264, -263, -263, -264,
  -263, -262, -262, -263,
  -262, -261, -261, -262,
  -261, -260, -260, -261,
  -280, -279, -279, -280,
  -279, -278, -278, -279,
  -278, -277, -277, -278,
  -277, -276, -276, -277,
  -276, -275, -275, -276,
  -275, -274, -274, -275,
  -274, -273, -273, -274,
  -273, -272, -272, -273,
  -272, -271, -271, -272,
  -271, -270, -270, -271,
  -270, -269, -269, -270,
  -269, -268, -268, -269,
  -268, -267, -267, -268,
  -267, -266, -266, -267,
  -266, -265, -265, -266,
  -265, -264, -264, -265,
  -264, -263, -263, -264,
  -263, -262, -262, -263,
  -262, -261, -261, -262,
  -261, -260, -260, -261,
  -280, -279, -279, -280,
  -279, -278, -278, -279,
  -278, -277, -277, -278,
  -277, -276, -276, -277,
  -276, -275, -275, -276,
  -275, -274, -274, -275,
  -274, -273, -273, -274,
  -273, -272, -272, -273,
  -272, -271, -271, -272,
  -271, -270, -270, -271,
  -270, -269, -269, -270,
  -269, -268, -268, -269,
  -268, -267, -267, -268,
  -267, -266, -266, -267,
  -266, -265, -265, -266,
  -265, -264, -264, -265,
  -264, -263, -263, -264,
  -263, -262, -262, -263,
  -262, -261, -261, -262,
  -261, -260, -260, -261,
  -280, -279, -279, -280,
  -279, -278, -278, -279,
  -278, -277, -277, -278,
  -277, -276, -276, -277,
  -276, -275, -275, -276,
  -275, -274, -274, -275,
  -274, -273, -273, -274,
  -273, -272, -272, -273,
  -272, -271, -271, -272,
  -271, -270, -270, -271,
  -270, -269, -269, -270,
  -269, -268, -268, -269,
  -268, -267, -267, -268,
  -267, -266, -266, -267,
  -266, -265, -265, -266,
  -265, -264, -264, -265,
  -264, -263, -263, -264,
  -263, -262, -262, -263,
  -262, -261, -261, -262,
  -261, -260, -260, -261,
  -280, -279, -279, -280,
  -279, -278, -278, -279,
  -278, -277, -277, -278,
  -277, -276, -276, -277,
  -276, -275, -275, -276,
  -275, -274, -274, -275,
  -274, -273, -273, -274,
  -273, -272, -272, -273,
  -272, -271, -271, -272,
  -271, -270, -270, -271,
  -270, -269, -269, -270,
  -269, -268, -268, -269,
  -268, -267, -267, -268,
  -267, -266, -266, -267,
  -266, -265, -265, -266,
  -265, -264, -264, -265,
  -264, -263, -263, -264,
  -263, -262, -262, -263,
  -262, -261, -261, -262,
  -261, -260, -260, -261,
  -280, -279, -279, -280,
  -279, -278, -278, -279,
  -278, -277, -277, -278,
  -277, -276, -276, -277,
  -276, -275, -275, -276,
  -275, -274, -274, -275,
  -274, -273, -273, -274,
  -273, -272, -272, -273,
  -272, -271, -271, -272,
  -271, -270, -270, -271,
  -270, -269, -269, -270,
  -269, -268, -268, -269,
  -268, -267, -267, -268,
  -267, -266, -266, -267,
  -266, -265, -265, -266,
  -265, -264, -264, -265,
  -264, -263, -263, -264,
  -263, -262, -262, -263,
  -262, -261, -261, -262,
  -261, -260, -260, -261,
  -280, -279, -279, -280,
  -279, -278, -278, -279,
  -278, -277, -277, -278,
  -277, -276, -276, -277,
  -276, -275, -275, -276,
  -275, -274, -274, -275,
  -274, -273, -273, -274,
  -273, -272, -272, -273,
  -272, -271, -271, -272,
  -271, -270, -270, -271,
  -270, -269, -269, -270,
  -269, -268, -268, -269,
  -268, -267, -267, -268,
  -267, -266, -266, -267,
  -266, -265, -265, -266,
  -265, -264, -264, -265,
  -264, -263, -263, -264,
  -263, -262, -262, -263,
  -262, -261, -261, -262,
  -261, -260, -260, -261 ;

 lat =
  -81.5, -81.5, -81.5, -81.5, -81.5, -81.5, -81.5, -81.5, -81.5, -81.5, 
    -81.5, -81.5, -81.5, -81.5, -81.5, -81.5, -81.5, -81.5, -81.5, -81.5,
  -80.5, -80.5, -80.5, -80.5, -80.5, -80.5, -80.5, -80.5, -80.5, -80.5, 
    -80.5, -80.5, -80.5, -80.5, -80.5, -80.5, -80.5, -80.5, -80.5, -80.5,
  -79.5, -79.5, -79.5, -79.5, -79.5, -79.5, -79.5, -79.5, -79.5, -79.5, 
    -79.5, -79.5, -79.5, -79.5, -79.5, -79.5, -79.5, -79.5, -79.5, -79.5,
  -78.5, -78.5, -78.5, -78.5, -78.5, -78.5, -78.5, -78.5, -78.5, -78.5, 
    -78.5, -78.5, -78.5, -78.5, -78.5, -78.5, -78.5, -78.5, -78.5, -78.5,
  -77.5, -77.5, -77.5, -77.5, -77.5, -77.5, -77.5, -77.5, -77.5, -77.5, 
    -77.5, -77.5, -77.5, -77.5, -77.5, -77.5, -77.5, -77.5, -77.5, -77.5,
  -76.5, -76.5, -76.5, -76.5, -76.5, -76.5, -76.5, -76.5, -76.5, -76.5, 
    -76.5, -76.5, -76.5, -76.5, -76.5, -76.5, -76.5, -76.5, -76.5, -76.5,
  -75.5, -75.5, -75.5, -75.5, -75.5, -75.5, -75.5, -75.5, -75.5, -75.5, 
    -75.5, -75.5, -75.5, -75.5, -75.5, -75.5, -75.5, -75.5, -75.5, -75.5,
  -74.5, -74.5, -74.5, -74.5, -74.5, -74.5, -74.5, -74.5, -74.5, -74.5, 
    -74.5, -74.5, -74.5, -74.5, -74.5, -74.5, -74.5, -74.5, -74.5, -74.5,
  -73.5, -73.5, -73.5, -73.5, -73.5, -73.5, -73.5, -73.5, -73.5, -73.5, 
    -73.5, -73.5, -73.5, -73.5, -73.5, -73.5, -73.5, -73.5, -73.5, -73.5,
  -72.5, -72.5, -72.5, -72.5, -72.5, -72.5, -72.5, -72.5, -72.5, -72.5, 
    -72.5, -72.5, -72.5, -72.5, -72.5, -72.5, -72.5, -72.5, -72.5, -72.5,
  -71.5, -71.5, -71.5, -71.5, -71.5, -71.5, -71.5, -71.5, -71.5, -71.5, 
    -71.5, -71.5, -71.5, -71.5, -71.5, -71.5, -71.5, -71.5, -71.5, -71.5,
  -70.5, -70.5, -70.5, -70.5, -70.5, -70.5, -70.5, -70.5, -70.5, -70.5, 
    -70.5, -70.5, -70.5, -70.5, -70.5, -70.5, -70.5, -70.5, -70.5, -70.5,
  -69.5, -69.5, -69.5, -69.5, -69.5, -69.5, -69.5, -69.5, -69.5, -69.5, 
    -69.5, -69.5, -69.5, -69.5, -69.5, -69.5, -69.5, -69.5, -69.5, -69.5,
  -68.5, -68.5, -68.5, -68.5, -68.5, -68.5, -68.5, -68.5, -68.5, -68.5, 
    -68.5, -68.5, -68.5, -68.5, -68.5, -68.5, -68.5, -68.5, -68.5, -68.5,
  -67.5, -67.5, -67.5, -67.5, -67.5, -67.5, -67.5, -67.5, -67.5, -67.5, 
    -67.5, -67.5, -67.5, -67.5, -67.5, -67.5, -67.5, -67.5, -67.5, -67.5,
  -66.5, -66.5, -66.5, -66.5, -66.5, -66.5, -66.5, -66.5, -66.5, -66.5, 
    -66.5, -66.5, -66.5, -66.5, -66.5, -66.5, -66.5, -66.5, -66.5, -66.5,
  -65.5, -65.5, -65.5, -65.5, -65.5, -65.5, -65.5, -65.5, -65.5, -65.5, 
    -65.5, -65.5, -65.5, -65.5, -65.5, -65.5, -65.5, -65.5, -65.5, -65.5,
  -64.5, -64.5, -64.5, -64.5, -64.5, -64.5, -64.5, -64.5, -64.5, -64.5, 
    -64.5, -64.5, -64.5, -64.5, -64.5, -64.5, -64.5, -64.5, -64.5, -64.5,
  -63.5, -63.5, -63.5, -63.5, -63.5, -63.5, -63.5, -63.5, -63.5, -63.5, 
    -63.5, -63.5, -63.5, -63.5, -63.5, -63.5, -63.5, -63.5, -63.5, -63.5,
  -62.5, -62.5, -62.5, -62.5, -62.5, -62.5, -62.5, -62.5, -62.5, -62.5, 
    -62.5, -62.5, -62.5, -62.5, -62.5, -62.5, -62.5, -62.5, -62.5, -62.5 ;

 lat_bnds =
  -82, -82, -81, -81,
  -82, -82, -81, -81,
  -82, -82, -81, -81,
  -82, -82, -81, -81,
  -82, -82, -81, -81,
  -82, -82, -81, -81,
  -82, -82, -81, -81,
  -82, -82, -81, -81,
  -82, -82, -81, -81,
  -82, -82, -81, -81,
  -82, -82, -81, -81,
  -82, -82, -81, -81,
  -82, -82, -81, -81,
  -82, -82, -81, -81,
  -82, -82, -81, -81,
  -82, -82, -81, -81,
  -82, -82, -81, -81,
  -82, -82, -81, -81,
  -82, -82, -81, -81,
  -82, -82, -81, -81,
  -81, -81, -80, -80,
  -81, -81, -80, -80,
  -81, -81, -80, -80,
  -81, -81, -80, -80,
  -81, -81, -80, -80,
  -81, -81, -80, -80,
  -81, -81, -80, -80,
  -81, -81, -80, -80,
  -81, -81, -80, -80,
  -81, -81, -80, -80,
  -81, -81, -80, -80,
  -81, -81, -80, -80,
  -81, -81, -80, -80,
  -81, -81, -80, -80,
  -81, -81, -80, -80,
  -81, -81, -80, -80,
  -81, -81, -80, -80,
  -81, -81, -80, -80,
  -81, -81, -80, -80,
  -81, -81, -80, -80,
  -80, -80, -79, -79,
  -80, -80, -79, -79,
  -80, -80, -79, -79,
  -80, -80, -79, -79,
  -80, -80, -79, -79,
  -80, -80, -79, -79,
  -80, -80, -79, -79,
  -80, -80, -79, -79,
  -80, -80, -79, -79,
  -80, -80, -79, -79,
  -80, -80, -79, -79,
  -80, -80, -79, -79,
  -80, -80, -79, -79,
  -80, -80, -79, -79,
  -80, -80, -79, -79,
  -80, -80, -79, -79,
  -80, -80, -79, -79,
  -80, -80, -79, -79,
  -80, -80, -79, -79,
  -80, -80, -79, -79,
  -79, -79, -78, -78,
  -79, -79, -78, -78,
  -79, -79, -78, -78,
  -79, -79, -78, -78,
  -79, -79, -78, -78,
  -79, -79, -78, -78,
  -79, -79, -78, -78,
  -79, -79, -78, -78,
  -79, -79, -78, -78,
  -79, -79, -78, -78,
  -79, -79, -78, -78,
  -79, -79, -78, -78,
  -79, -79, -78, -78,
  -79, -79, -78, -78,
  -79, -79, -78, -78,
  -79, -79, -78, -78,
  -79, -79, -78, -78,
  -79, -79, -78, -78,
  -79, -79, -78, -78,
  -79, -79, -78, -78,
  -78, -78, -77, -77,
  -78, -78, -77, -77,
  -78, -78, -77, -77,
  -78, -78, -77, -77,
  -78, -78, -77, -77,
  -78, -78, -77, -77,
  -78, -78, -77, -77,
  -78, -78, -77, -77,
  -78, -78, -77, -77,
  -78, -78, -77, -77,
  -78, -78, -77, -77,
  -78, -78, -77, -77,
  -78, -78, -77, -77,
  -78, -78, -77, -77,
  -78, -78, -77, -77,
  -78, -78, -77, -77,
  -78, -78, -77, -77,
  -78, -78, -77, -77,
  -78, -78, -77, -77,
  -78, -78, -77, -77,
  -77, -77, -76, -76,
  -77, -77, -76, -76,
  -77, -77, -76, -76,
  -77, -77, -76, -76,
  -77, -77, -76, -76,
  -77, -77, -76, -76,
  -77, -77, -76, -76,
  -77, -77, -76, -76,
  -77, -77, -76, -76,
  -77, -77, -76, -76,
  -77, -77, -76, -76,
  -77, -77, -76, -76,
  -77, -77, -76, -76,
  -77, -77, -76, -76,
  -77, -77, -76, -76,
  -77, -77, -76, -76,
  -77, -77, -76, -76,
  -77, -77, -76, -76,
  -77, -77, -76, -76,
  -77, -77, -76, -76,
  -76, -76, -75, -75,
  -76, -76, -75, -75,
  -76, -76, -75, -75,
  -76, -76, -75, -75,
  -76, -76, -75, -75,
  -76, -76, -75, -75,
  -76, -76, -75, -75,
  -76, -76, -75, -75,
  -76, -76, -75, -75,
  -76, -76, -75, -75,
  -76, -76, -75, -75,
  -76, -76, -75, -75,
  -76, -76, -75, -75,
  -76, -76, -75, -75,
  -76, -76, -75, -75,
  -76, -76, -75, -75,
  -76, -76, -75, -75,
  -76, -76, -75, -75,
  -76, -76, -75, -75,
  -76, -76, -75, -75,
  -75, -75, -74, -74,
  -75, -75, -74, -74,
  -75, -75, -74, -74,
  -75, -75, -74, -74,
  -75, -75, -74, -74,
  -75, -75, -74, -74,
  -75, -75, -74, -74,
  -75, -75, -74, -74,
  -75, -75, -74, -74,
  -75, -75, -74, -74,
  -75, -75, -74, -74,
  -75, -75, -74, -74,
  -75, -75, -74, -74,
  -75, -75, -74, -74,
  -75, -75, -74, -74,
  -75, -75, -74, -74,
  -75, -75, -74, -74,
  -75, -75, -74, -74,
  -75, -75, -74, -74,
  -75, -75, -74, -74,
  -74, -74, -73, -73,
  -74, -74, -73, -73,
  -74, -74, -73, -73,
  -74, -74, -73, -73,
  -74, -74, -73, -73,
  -74, -74, -73, -73,
  -74, -74, -73, -73,
  -74, -74, -73, -73,
  -74, -74, -73, -73,
  -74, -74, -73, -73,
  -74, -74, -73, -73,
  -74, -74, -73, -73,
  -74, -74, -73, -73,
  -74, -74, -73, -73,
  -74, -74, -73, -73,
  -74, -74, -73, -73,
  -74, -74, -73, -73,
  -74, -74, -73, -73,
  -74, -74, -73, -73,
  -74, -74, -73, -73,
  -73, -73, -72, -72,
  -73, -73, -72, -72,
  -73, -73, -72, -72,
  -73, -73, -72, -72,
  -73, -73, -72, -72,
  -73, -73, -72, -72,
  -73, -73, -72, -72,
  -73, -73, -72, -72,
  -73, -73, -72, -72,
  -73, -73, -72, -72,
  -73, -73, -72, -72,
  -73, -73, -72, -72,
  -73, -73, -72, -72,
  -73, -73, -72, -72,
  -73, -73, -72, -72,
  -73, -73, -72, -72,
  -73, -73, -72, -72,
  -73, -73, -72, -72,
  -73, -73, -72, -72,
  -73, -73, -72, -72,
  -72, -72, -71, -71,
  -72, -72, -71, -71,
  -72, -72, -71, -71,
  -72, -72, -71, -71,
  -72, -72, -71, -71,
  -72, -72, -71, -71,
  -72, -72, -71, -71,
  -72, -72, -71, -71,
  -72, -72, -71, -71,
  -72, -72, -71, -71,
  -72, -72, -71, -71,
  -72, -72, -71, -71,
  -72, -72, -71, -71,
  -72, -72, -71, -71,
  -72, -72, -71, -71,
  -72, -72, -71, -71,
  -72, -72, -71, -71,
  -72, -72, -71, -71,
  -72, -72, -71, -71,
  -72, -72, -71, -71,
  -71, -71, -70, -70,
  -71, -71, -70, -70,
  -71, -71, -70, -70,
  -71, -71, -70, -70,
  -71, -71, -70, -70,
  -71, -71, -70, -70,
  -71, -71, -70, -70,
  -71, -71, -70, -70,
  -71, -71, -70, -70,
  -71, -71, -70, -70,
  -71, -71, -70, -70,
  -71, -71, -70, -70,
  -71, -71, -70, -70,
  -71, -71, -70, -70,
  -71, -71, -70, -70,
  -71, -71, -70, -70,
  -71, -71, -70, -70,
  -71, -71, -70, -70,
  -71, -71, -70, -70,
  -71, -71, -70, -70,
  -70, -70, -69, -69,
  -70, -70, -69, -69,
  -70, -70, -69, -69,
  -70, -70, -69, -69,
  -70, -70, -69, -69,
  -70, -70, -69, -69,
  -70, -70, -69, -69,
  -70, -70, -69, -69,
  -70, -70, -69, -69,
  -70, -70, -69, -69,
  -70, -70, -69, -69,
  -70, -70, -69, -69,
  -70, -70, -69, -69,
  -70, -70, -69, -69,
  -70, -70, -69, -69,
  -70, -70, -69, -69,
  -70, -70, -69, -69,
  -70, -70, -69, -69,
  -70, -70, -69, -69,
  -70, -70, -69, -69,
  -69, -69, -68, -68,
  -69, -69, -68, -68,
  -69, -69, -68, -68,
  -69, -69, -68, -68,
  -69, -69, -68, -68,
  -69, -69, -68, -68,
  -69, -69, -68, -68,
  -69, -69, -68, -68,
  -69, -69, -68, -68,
  -69, -69, -68, -68,
  -69, -69, -68, -68,
  -69, -69, -68, -68,
  -69, -69, -68, -68,
  -69, -69, -68, -68,
  -69, -69, -68, -68,
  -69, -69, -68, -68,
  -69, -69, -68, -68,
  -69, -69, -68, -68,
  -69, -69, -68, -68,
  -69, -69, -68, -68,
  -68, -68, -67, -67,
  -68, -68, -67, -67,
  -68, -68, -67, -67,
  -68, -68, -67, -67,
  -68, -68, -67, -67,
  -68, -68, -67, -67,
  -68, -68, -67, -67,
  -68, -68, -67, -67,
  -68, -68, -67, -67,
  -68, -68, -67, -67,
  -68, -68, -67, -67,
  -68, -68, -67, -67,
  -68, -68, -67, -67,
  -68, -68, -67, -67,
  -68, -68, -67, -67,
  -68, -68, -67, -67,
  -68, -68, -67, -67,
  -68, -68, -67, -67,
  -68, -68, -67, -67,
  -68, -68, -67, -67,
  -67, -67, -66, -66,
  -67, -67, -66, -66,
  -67, -67, -66, -66,
  -67, -67, -66, -66,
  -67, -67, -66, -66,
  -67, -67, -66, -66,
  -67, -67, -66, -66,
  -67, -67, -66, -66,
  -67, -67, -66, -66,
  -67, -67, -66, -66,
  -67, -67, -66, -66,
  -67, -67, -66, -66,
  -67, -67, -66, -66,
  -67, -67, -66, -66,
  -67, -67, -66, -66,
  -67, -67, -66, -66,
  -67, -67, -66, -66,
  -67, -67, -66, -66,
  -67, -67, -66, -66,
  -67, -67, -66, -66,
  -66, -66, -65, -65,
  -66, -66, -65, -65,
  -66, -66, -65, -65,
  -66, -66, -65, -65,
  -66, -66, -65, -65,
  -66, -66, -65, -65,
  -66, -66, -65, -65,
  -66, -66, -65, -65,
  -66, -66, -65, -65,
  -66, -66, -65, -65,
  -66, -66, -65, -65,
  -66, -66, -65, -65,
  -66, -66, -65, -65,
  -66, -66, -65, -65,
  -66, -66, -65, -65,
  -66, -66, -65, -65,
  -66, -66, -65, -65,
  -66, -66, -65, -65,
  -66, -66, -65, -65,
  -66, -66, -65, -65,
  -65, -65, -64, -64,
  -65, -65, -64, -64,
  -65, -65, -64, -64,
  -65, -65, -64, -64,
  -65, -65, -64, -64,
  -65, -65, -64, -64,
  -65, -65, -64, -64,
  -65, -65, -64, -64,
  -65, -65, -64, -64,
  -65, -65, -64, -64,
  -65, -65, -64, -64,
  -65, -65, -64, -64,
  -65, -65, -64, -64,
  -65, -65, -64, -64,
  -65, -65, -64, -64,
  -65, -65, -64, -64,
  -65, -65, -64, -64,
  -65, -65, -64, -64,
  -65, -65, -64, -64,
  -65, -65, -64, -64,
  -64, -64, -63, -63,
  -64, -64, -63, -63,
  -64, -64, -63, -63,
  -64, -64, -63, -63,
  -64, -64, -63, -63,
  -64, -64, -63, -63,
  -64, -64, -63, -63,
  -64, -64, -63, -63,
  -64, -64, -63, -63,
  -64, -64, -63, -63,
  -64, -64, -63, -63,
  -64, -64, -63, -63,
  -64, -64, -63, -63,
  -64, -64, -63, -63,
  -64, -64, -63, -63,
  -64, -64, -63, -63,
  -64, -64, -63, -63,
  -64, -64, -63, -63,
  -64, -64, -63, -63,
  -64, -64, -63, -63,
  -63, -63, -62, -62,
  -63, -63, -62, -62,
  -63, -63, -62, -62,
  -63, -63, -62, -62,
  -63, -63, -62, -62,
  -63, -63, -62, -62,
  -63, -63, -62, -62,
  -63, -63, -62, -62,
  -63, -63, -62, -62,
  -63, -63, -62, -62,
  -63, -63, -62, -62,
  -63, -63, -62, -62,
  -63, -63, -62, -62,
  -63, -63, -62, -62,
  -63, -63, -62, -62,
  -63, -63, -62, -62,
  -63, -63, -62, -62,
  -63, -63, -62, -62,
  -63, -63, -62, -62,
  -63, -63, -62, -62 ;

 time = 49290.5, 49320, 49349.5, 49380 ;

 time_bnds =
  49275, 49306,
  49306, 49334,
  49334, 49365,
  49365, 49395 ;

 average_DT = 31, 28, 31, 30 ;

 zsatcalc =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  50.03294, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  53.57268, 53.30359, 53.11386, 52.48583, 49.4257, _, _, _, _, 45.92426, 
    55.98218, 52.89568, 52.72888, 48.16253, _, _, _, _, _, _,
  39.9788, 40.10589, 43.3566, 44.80859, 49.80643, 52.41396, 53.16078, 
    55.38807, 55.44016, 54.54989, 49.93708, 48.50716, 49.83224, 49.79397, 
    51.41099, _, _, _, _, _,
  39.98369, 39.98371, 39.98296, 39.98288, 39.98311, 42.6967, 46.48512, 
    47.80087, 48.15093, 47.29153, 46.6727, 44.84358, 48.20004, 49.51279, 
    53.66824, 54.40544, 53.27378, 53.15202, 54.48359, 55.45014,
  39.98312, 40.46659, 39.98295, 39.98299, 39.98284, 39.98301, 42.42885, 
    43.87981, 46.11009, 45.94758, 47.60431, 46.69874, 48.02461, 46.13491, 
    45.21923, 44.35905, 43.38848, 39.97417, 41.12476, 46.27187,
  39.21393, 39.28007, 39.5602, 39.21997, 39.7663, 39.98232, 40.81654, 
    39.84905, 39.71074, 38.46192, 37.49322, 38.57851, 41.26633, 46.3688, 
    47.26487, 47.72254, 48.153, 48.5554, 48.4213, 48.55573,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  59.71378, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  58.73066, 59.003, 59.53012, 58.61917, 49.42974, _, _, _, _, 59.53199, 
    69.30826, 59.27387, 59.16808, 48.63815, _, _, _, _, _, _,
  39.94944, 39.97241, 43.98794, 49.96777, 59.16006, 58.86485, 57.69952, 
    57.72708, 57.54683, 57.66161, 49.94027, 49.90716, 49.84163, 59.5921, 
    59.67007, _, _, _, _, _,
  39.98372, 39.98377, 39.98312, 39.98317, 39.98352, 39.98328, 43.22574, 
    43.6414, 43.25522, 40.19134, 39.98235, 39.98065, 49.97383, 49.97046, 
    59.1527, 59.31867, 59.40725, 59.7867, 59.77913, 59.45736,
  39.95356, 39.98313, 39.98317, 39.9832, 39.98303, 39.98316, 39.9837, 
    39.98356, 39.98353, 39.98396, 41.35232, 41.5306, 41.85748, 39.98187, 
    39.9801, 39.97982, 39.9769, 39.97471, 39.97047, 45.04634,
  39.92108, 39.77235, 39.98064, 39.95094, 39.98141, 39.98238, 39.98353, 
    39.98332, 39.9832, 39.98434, 39.98383, 39.98402, 43.49437, 48.19402, 
    49.44313, 49.97957, 49.98013, 49.97944, 49.9797, 49.89053,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  59.95761, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  49.8055, 49.33381, 49.15622, 48.99057, 48.7038, _, _, _, _, 58.85986, 
    58.67538, 58.58006, 58.6368, 47.98195, _, _, _, _, _, _,
  39.73877, 36.04705, 39.72803, 46.76117, 49.40855, 49.45325, 49.54664, 
    49.2803, 49.54982, 51.40908, 46.38293, 48.63297, 51.02205, 57.34545, 
    59.69253, _, _, _, _, _,
  30.64117, 29.93299, 31.8317, 37.32819, 39.9224, 39.74264, 39.52189, 
    37.46815, 41.19892, 42.37855, 43.76529, 43.40236, 46.965, 49.97115, 
    49.96427, 53.52724, 53.34009, 54.67731, 56.57291, 57.41077,
  29.30867, 31.15795, 29.36013, 30.96096, 36.97813, 39.21212, 39.98368, 
    39.98351, 39.98343, 39.98384, 39.9837, 39.98351, 41.72979, 42.58821, 
    43.25816, 41.88768, 41.88473, 42.15118, 43.54367, 47.10654,
  34.75978, 32.51633, 34.58174, 35.19574, 36.25374, 39.29942, 39.51448, 
    38.89968, 39.98309, 39.9842, 39.98367, 40.68251, 44.95482, 47.18433, 
    49.468, 49.97953, 49.98013, 49.97946, 49.97973, 49.9798,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  56.84623, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, 54.50643, 56.44537, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, 38.37991, 46.71422, 50.06669, 51.73561, 
    48.6559, 49.47305, 56.30112, 57.67973,
  _, _, _, _, _, _, 29.98753, 37.48435, 29.98755, 30.21004, 30.59978, 
    35.41387, 41.14043, 44.23502, 45.03118, 42.50593, 36.10816, 40.40921, 
    44.80895, 47.60775,
  _, _, _, _, _, _, _, 19.99151, 23.87872, 31.65411, 38.66061, 39.35899, 
    39.3172, 42.27552, 43.1559, 47.69215, 46.73336, 46.52934, 46.42954, 
    45.48595 ;
}
