netcdf tas_daily_exAA06_senC2CH4rcp85_r1i1p1_20010101-20501231_box {
dimensions:
	lon = 20 ;
	bnds = 2 ;
	lat = 20 ;
	time = UNLIMITED ; // (4 currently)
variables:
	double lon(lon) ;
		lon:standard_name = "longitude" ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:axis = "X" ;
		lon:bounds = "lon_bnds" ;
	double lon_bnds(lon, bnds) ;
	double lat(lat) ;
		lat:standard_name = "latitude" ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:axis = "Y" ;
		lat:bounds = "lat_bnds" ;
	double lat_bnds(lat, bnds) ;
	double height ;
		height:standard_name = "height" ;
		height:long_name = "height" ;
		height:units = "m" ;
		height:positive = "up" ;
		height:axis = "Z" ;
	double time(time) ;
		time:standard_name = "time" ;
		time:long_name = "time" ;
		time:bounds = "time_bnds" ;
		time:units = "days since 1860-1-1 00:00:00" ;
		time:calendar = "365_day" ;
		time:axis = "T" ;
	double time_bnds(time, bnds) ;
	float tas(time, lat, lon) ;
		tas:standard_name = "air_temperature" ;
		tas:long_name = "Near-Surface Air Temperature" ;
		tas:units = "K" ;
		tas:grid_type = "gaussian" ;
		tas:coordinates = "height" ;
		tas:_FillValue = 1.e+20f ;
		tas:missing_value = 1.e+20f ;
		tas:comment = "near-surface (usually, 2 meter) air temperature" ;
		tas:cell_methods = "time: point" ;
		tas:history = "2017-03-14T00:18:28Z altered by CMOR: Treated scalar dimension: \'height\'. 2017-03-14T00:18:28Z altered by CMOR: replaced missing value flag (1e+38) with standard missing value (1e+20)." ;
		tas:associated_files = "baseURL: http://www.met.reading.ac.uk/ccmi/ gridspecFile: gridspec_atmos_fx_CMAM_senC2CH4rcp85_r0i0p0.nc areacella: areacella_fx_CMAM_senC2CH4rcp85_r0i0p0.nc" ;

// global attributes:
		:CDI = "Climate Data Interface version ?? (http://mpimet.mpg.de/cdi)" ;
		:Conventions = "CF-1.4" ;
		:history = "reset by cdo to create anonymous sample file" ;
		:source = "201707_compliance_checker_evaluation/work/p1.py" ;
		:institution = "CEDA" ;
		:institute_id = "CEDA" ;
		:experiment_id = "senC2CH4rcp85" ;
		:model_id = "exAA06" ;
		:forcing = "N/A" ;
		:parent_experiment_id = "N/A" ;
		:parent_experiment_rip = "N/A" ;
		:branch_time = 0. ;
		:contact = "none" ;
		:references = "http://www.cccma.ec.gc.ca/models" ;
		:initialization_method = 1 ;
		:physics_version = 1 ;
		:tracking_id = "3ddea2ef-56a6-4642-b985-e6f3cef49563" ;
		:CCCma_runid = "ccmi1_dp962q" ;
		:CCCma_data_licence = "1) GRANT OF LICENCE - The Government of Canada (Environment Canada) is the \n",
			"owner of all intellectual property rights (including copyright) that may exist in this Data \n",
			"product. You (as \"The Licensee\") are hereby granted a non-exclusive, non-assignable, \n",
			"non-transferable unrestricted licence to use this data product for any purpose including \n",
			"the right to share these data with others and to make value-added and derivative \n",
			"products from it. This licence is not a sale of any or all of the owner\'s rights.\n",
			"2) NO WARRANTY - This Data product is provided \"as-is\"; it has not been designed or \n",
			"prepared to meet the Licensee\'s particular requirements. Environment Canada makes no \n",
			"warranty, either express or implied, including but not limited to, warranties of \n",
			"merchantability and fitness for a particular purpose. In no event will Environment Canada \n",
			"be liable for any indirect, special, consequential or other damages attributed to the \n",
			"Licensee\'s use of the Data product." ;
		:product = "output" ;
		:experiment = "Projection Scenario - CH4-RCP8.5" ;
		:frequency = "day" ;
		:creation_date = "2017-03-14T00:18:28Z" ;
		:project_id = "CCMI1" ;
		:table_id = "Table daily (31 October 2014) cb63dd622146f1647dc224701f367b1c" ;
		:title = "Dummy file with known metadata errors" ;
		:parent_experiment = "N/A" ;
		:modeling_realm = "atmos" ;
		:realization = 1 ;
		:cmor_version = "2.8.2" ;
		:comment = "this is a sample file with known metadata errors" ;
		:CDO = "Climate Data Operators version 1.7.0 (http://mpimet.mpg.de/cdo)" ;
data:

 lon = 0, 3.75, 7.5, 11.25, 15, 18.75, 22.5, 26.25, 30, 33.75, 37.5, 41.25, 
    45, 48.75, 52.5, 56.25, 60, 63.75, 67.5, 71.25 ;

 lon_bnds =
  0, 1.875,
  1.875, 5.625,
  5.625, 9.375,
  9.375, 13.125,
  13.125, 16.875,
  16.875, 20.625,
  20.625, 24.375,
  24.375, 28.125,
  28.125, 31.875,
  31.875, 35.625,
  35.625, 39.375,
  39.375, 43.125,
  43.125, 46.875,
  46.875, 50.625,
  50.625, 54.375,
  54.375, 58.125,
  58.125, 61.875,
  61.875, 65.625,
  65.625, 69.375,
  69.375, 73.125 ;

 lat = -87.1590944530229, -83.4789365664772, -79.7770455519856, 
    -76.0702443597051, -72.3615809265049, -68.6520166866775, 
    -64.9419493859175, -61.2315730852371, -57.52099369513, -53.8102739291014, 
    -50.0994533101468, -46.3885580087654, -42.6776060697649, 
    -38.966610366614, -35.2555803585282, -31.5445231811817, 
    -27.8334443491532, -24.122348223248, -20.4112383307278, -16.7001175910027 ;

 lat_bnds =
  -90, -85.31901550975,
  -85.31901550975, -81.6279910592314,
  -81.6279910592314, -77.9236449558454,
  -77.9236449558454, -74.215912643105,
  -74.215912643105, -70.5067988065912,
  -70.5067988065912, -66.7969830362975,
  -66.7969830362975, -63.0867612355773,
  -63.0867612355773, -59.3762833901836,
  -59.3762833901836, -55.6656338121157,
  -55.6656338121157, -51.9548636196241,
  -51.9548636196241, -48.2440056594561,
  -48.2440056594561, -44.5330820392652,
  -44.5330820392652, -40.8221082181895,
  -40.8221082181895, -37.1110953625711,
  -37.1110953625711, -33.4000517698549,
  -33.4000517698549, -29.6889837651674,
  -29.6889837651674, -25.9778962862006,
  -25.9778962862006, -22.2667932769879,
  -22.2667932769879, -18.5556779608652,
  -18.5556779608652, -14.8445530351254 ;

 height = 2 ;

 time = 51465, 51466, 51467, 51468 ;

 time_bnds =
  51464.5, 51465.5,
  51465.5, 51466.5,
  51466.5, 51467.5,
  51467.5, 51468.5 ;

 tas =
  251.7849, 251.4744, 251.1742, 250.8769, 250.5958, 250.3883, 250.1382, 
    249.9572, 249.7202, 249.576, 249.3612, 249.2317, 249.008, 248.9006, 
    248.7372, 248.6327, 248.5695, 248.568, 248.8461, 249.1861,
  250.0131, 249.3097, 248.5827, 248.078, 247.4717, 246.8345, 246.0781, 
    245.0215, 243.7177, 242.7611, 242.2137, 242.0327, 241.9591, 242.1637, 
    242.1254, 242.0709, 242.2255, 242.1754, 242.3255, 242.3388,
  248.1868, 247.6291, 247.3569, 246.6137, 245.5321, 243.2202, 240.8672, 
    239.1807, 239.0218, 240.305, 242.2063, 243.6249, 244.6845, 246.6947, 
    247.9028, 248.465, 248.4591, 248.0794, 247.4334, 246.7359,
  246.5813, 246.6167, 245.6278, 243.9354, 240.7583, 237.3486, 231.6977, 
    235.0132, 239.2411, 243.2364, 244.8434, 245.8338, 245.9177, 245.2481, 
    245.5218, 246.7771, 249.0124, 251.0211, 251.7746, 251.2124,
  252.3043, 252.3397, 252.556, 254.2101, 254.7428, 254.5809, 254.4587, 
    254.2704, 253.5905, 253.4316, 253.0048, 250.9976, 246.2914, 243.1025, 
    246.6255, 250.8063, 250.5988, 249.9925, 253.1343, 255.0842,
  270.2533, 270.3533, 263.9299, 263.6414, 264.0005, 264.0388, 263.8327, 
    263.6444, 263.2971, 262.4671, 261.047, 259.4533, 257.8051, 255.4697, 
    252.5163, 251.7113, 254.859, 258.897, 261.3193, 262.2419,
  272.1825, 272.3238, 271.7675, 272.415, 270.6079, 270.577, 272.2958, 
    272.0986, 269.1849, 269.0363, 269.3423, 269.722, 269.8088, 269.338, 
    268.4315, 267.444, 266.7671, 266.7082, 266.5346, 266.1328,
  273.8954, 274.3148, 274.2251, 273.9602, 273.8469, 273.9602, 274.2413, 
    274.1809, 273.8351, 273.5452, 273.476, 273.5526, 273.607, 272.9242, 
    272.4312, 271.6425, 271.1495, 270.7227, 270.4755, 270.3342,
  274.5665, 274.8578, 275.0874, 275.1066, 274.8402, 274.5782, 274.721, 
    275.2876, 275.7335, 275.8217, 275.6584, 275.6805, 275.9395, 275.9895, 
    275.7305, 275.4921, 275.5068, 275.5451, 275.5083, 275.6157,
  274.5415, 274.696, 275.2199, 275.548, 275.4274, 275.1272, 275.3965, 
    276.0101, 276.5281, 276.5752, 276.2882, 276.1735, 276.5384, 277.2109, 
    277.2374, 276.8754, 276.7386, 276.7459, 276.7915, 276.9799,
  276.0116, 276.4207, 276.6355, 276.7253, 276.9343, 277.1918, 277.9173, 
    278.0203, 279.5184, 279.6228, 278.8076, 277.9791, 277.5744, 277.6436, 
    278.0556, 278.1086, 277.8569, 278.0586, 278.6045, 279.2549,
  278.319, 278.6104, 278.681, 278.4927, 278.5118, 278.8988, 279.7155, 
    279.9348, 280.3557, 281.1724, 281.7125, 281.2651, 279.6817, 278.7473, 
    278.6487, 278.9547, 278.6428, 278.6384, 280.1644, 281.8288,
  282.1451, 282.0024, 281.8376, 281.6816, 281.7699, 282.3571, 283.1532, 
    283.5785, 284.2348, 284.7248, 285.3826, 285.7446, 284.7322, 283.4034, 
    282.7779, 282.4777, 282.179, 282.3997, 283.8684, 284.9603,
  285.6299, 285.4003, 285.3606, 285.518, 286.373, 288.3008, 290.3507, 
    291.475, 291.7487, 291.706, 291.3749, 291.4735, 290.7966, 289.9269, 
    289.3839, 288.0653, 287.54, 287.743, 289.0645, 289.0263,
  287.696, 287.9506, 288.2802, 288.9144, 290.002, 291.1262, 292.4197, 
    294.555, 296.7565, 296.4622, 293.8899, 293.004, 292.3771, 291.9341, 
    291.7487, 291.3646, 290.9614, 290.9864, 290.8805, 290.6141,
  291.0526, 291.1439, 291.188, 290.8658, 291.2999, 292.6567, 288.6098, 
    290.7686, 295.488, 298.518, 294.9774, 294.0885, 294.0444, 293.7074, 
    293.3792, 293.182, 293.2071, 292.8627, 292.6434, 292.4786,
  293.2379, 292.77, 291.5898, 290.7716, 291.5868, 292.3035, 291.4353, 
    288.9645, 292.6111, 298.9654, 298.0633, 297.2657, 297.2436, 297.304, 
    296.9125, 296.2017, 295.9825, 295.9516, 295.8191, 295.8073,
  293.4101, 292.9113, 291.9606, 292.3844, 294.3946, 292.1593, 293.3263, 
    290.9555, 291.2425, 295.5424, 300.2824, 300.3546, 296.1046, 298.4253, 
    299.3377, 298.5504, 298.3473, 298.5445, 298.3679, 298.3797,
  294.3446, 294.2122, 294.0503, 295.6896, 293.4307, 290.0755, 292.3197, 
    294.7125, 294.8714, 291.503, 300.7666, 301.4965, 293.5779, 293.575, 
    299.8189, 299.9352, 299.8056, 299.7379, 299.6011, 299.5584,
  296.1664, 296.1061, 296.627, 298.3149, 293.3145, 292.6993, 293.5426, 
    294.7007, 294.3976, 292.9466, 296.8227, 301.5936, 293.107, 294.9332, 
    300.0558, 300.381, 300.3634, 300.2883, 300.4944, 300.5959,
  248.2629, 247.9016, 247.5537, 247.2342, 246.924, 246.6274, 246.6018, 
    246.4467, 246.289, 246.0557, 245.8616, 245.9209, 245.7551, 245.6162, 
    245.7294, 245.6539, 245.8252, 245.7915, 246.0328, 246.1865,
  250.4796, 249.9753, 249.5142, 249.0342, 248.0984, 247.3326, 246.4791, 
    245.4234, 244.609, 243.7285, 242.8643, 241.5658, 239.8494, 238.7357, 
    239.8022, 241.4364, 242.871, 243.7973, 244.64, 245.0782,
  247.5321, 246.5775, 246.4333, 246.2324, 246.0139, 245.9384, 245.5488, 
    244.458, 245.1038, 245.3411, 245.027, 244.6117, 243.9443, 243.1097, 
    240.5802, 240.347, 242.5434, 243.9685, 245.0405, 245.8238,
  241.8921, 236.3371, 237.0652, 239.3074, 239.7321, 238.9663, 238.853, 
    239.9088, 241.1007, 242.1577, 243.022, 244.1721, 245.6243, 246.0544, 
    245.4234, 246.2526, 247.9771, 249.3699, 250.2328, 251.2818,
  252.622, 252.3402, 252.5533, 252.9686, 252.9645, 252.293, 251.6796, 
    251.8791, 252.5371, 253.2571, 253.1694, 251.8791, 249.8755, 250.7897, 
    250.1317, 247.8854, 248.6189, 250.0683, 251.4261, 252.1528,
  269.8225, 270.049, 260.3627, 260.7901, 261.347, 261.6706, 261.2944, 
    260.2886, 258.9052, 257.2184, 255.7757, 255.7326, 260.6796, 259.9785, 
    257.2346, 257.534, 258.8931, 259.3704, 261.1973, 262.6899,
  270.6693, 271.1263, 271.1317, 271.0994, 272.3816, 270.4576, 269.4275, 
    269.3668, 270.3929, 270.3564, 270.7218, 270.5722, 269.7834, 268.6751, 
    267.9605, 267.4468, 267.2337, 267.68, 268.4553, 269.4612,
  273.9699, 274.1776, 274.1223, 273.9672, 273.8095, 273.7218, 273.8419, 
    273.8351, 273.7003, 273.5519, 273.4468, 273.4144, 273.4899, 272.9695, 
    272.8522, 272.4234, 271.129, 270.8027, 271.0576, 271.454,
  275.1052, 275.1834, 275.1335, 275.0203, 274.9583, 275.0648, 275.3439, 
    275.6769, 275.7834, 275.6998, 275.5515, 275.596, 275.8818, 275.9884, 
    275.7726, 275.4477, 275.1753, 275.0499, 274.9461, 275.1457,
  274.903, 274.9879, 275.2185, 275.4383, 275.7416, 275.9911, 276.2513, 
    276.3295, 276.4239, 276.5317, 276.5398, 276.5452, 276.7677, 276.8769, 
    276.7906, 276.7664, 276.8257, 276.8135, 276.4279, 276.1529,
  276.3821, 276.7367, 276.7974, 276.8459, 277.0913, 277.1223, 276.978, 
    277.005, 277.4055, 277.7196, 277.5929, 277.5255, 278.1052, 278.5717, 
    278.6904, 278.5583, 278.6769, 278.658, 277.8908, 277.2328,
  278.6675, 278.863, 278.7618, 278.4881, 278.3843, 278.48, 278.5003, 
    278.5933, 278.9264, 279.2513, 279.4279, 279.5425, 280.0724, 280.3677, 
    280.0077, 279.9416, 280.9313, 282.0086, 281.9236, 281.0675,
  281.9317, 281.8967, 281.6108, 281.2306, 281.2077, 281.6769, 282.2473, 
    282.5385, 282.5627, 282.3133, 282.0949, 282.2499, 282.6747, 283.4001, 
    284.2967, 285.0612, 285.8001, 286.3947, 286.2962, 285.2742,
  285.3039, 285.1246, 285.1502, 285.285, 286.2841, 288.1043, 289.6387, 
    290.3088, 290.2873, 289.3434, 288.5399, 288.7515, 289.1345, 289.996, 
    290.6958, 290.6311, 290.0041, 289.307, 288.6342, 288.0234,
  287.9506, 287.8306, 288.072, 288.8769, 290.1915, 291.0194, 292.063, 
    293.7497, 294.9403, 294.1138, 293.2981, 293.143, 293.1053, 292.601, 
    292.3367, 291.7812, 291.0963, 290.8724, 290.3439, 289.8019,
  291.2459, 291.2648, 291.2041, 290.9318, 291.2271, 290.6028, 290.4437, 
    289.8383, 291.6518, 297.6086, 295.5012, 294.854, 294.4387, 294.0531, 
    293.9911, 293.6783, 293.0297, 292.7129, 292.5902, 292.4554,
  293.4059, 292.9987, 291.8931, 291.1313, 292.1493, 292.2652, 289.2599, 
    288.6733, 292.1938, 299.2711, 298.9124, 297.8635, 298.3313, 297.6639, 
    297.0248, 296.4235, 295.8666, 295.8154, 295.7142, 295.7938,
  293.6648, 292.7641, 291.8742, 292.4688, 293.9331, 291.8715, 292.3664, 
    290.8657, 292.9623, 298.9084, 300.3713, 300.2999, 297.0491, 298.5983, 
    299.081, 298.601, 298.5066, 298.5093, 298.179, 298.2558,
  294.4927, 293.9763, 293.9142, 295.899, 293.6136, 291.6963, 292.9165, 
    293.1727, 297.5898, 296.7713, 300.8594, 301.3327, 292.6468, 293.8199, 
    299.8199, 300.0167, 299.9587, 299.7255, 299.5151, 299.5583,
  296.3304, 296.0904, 296.5637, 298.2841, 293.147, 291.5951, 292.5187, 
    293.6904, 295.8949, 292.7102, 299.1349, 301.9124, 295.1911, 296.2697, 
    300.1596, 300.3673, 300.3713, 300.3902, 300.5641, 300.5978,
  251.0514, 250.5701, 249.8879, 249.3889, 248.6727, 248.1598, 247.4372, 
    246.8144, 246.2081, 245.7432, 245.1103, 244.7439, 244.4142, 244.1313, 
    244.1388, 243.9873, 244.1325, 244.226, 244.3953, 244.7604,
  251.3356, 249.994, 248.6234, 247.1744, 246.0148, 244.9145, 244.2892, 
    242.1707, 241.5984, 242.177, 243.4314, 243.5287, 243.7674, 244.0782, 
    243.6651, 243.9418, 243.9784, 243.9948, 243.9683, 243.7232,
  253.2065, 251.9533, 250.7406, 248.7535, 247.1997, 246.0981, 245.7267, 
    246.2017, 245.8253, 244.442, 242.5383, 240.9074, 239.4206, 237.6167, 
    238.0096, 240.2922, 242.5775, 245.2745, 246.3041, 246.7083,
  249.5039, 246.0767, 241.4595, 237.268, 231.4646, 237.8112, 242.4082, 
    245.2556, 245.6358, 245.4829, 243.6702, 241.3698, 240.9668, 242.4941, 
    244.677, 246.4582, 248.6019, 249.8361, 250.5271, 249.5759,
  253.7168, 252.4839, 252.0291, 251.0589, 249.4938, 249.7313, 251.1625, 
    252.0354, 252.9576, 253.2166, 249.9511, 247.2477, 248.5918, 249.9018, 
    249.8993, 250.09, 251.7487, 253.6145, 254.4331, 255.8884,
  270.014, 269.678, 257.5179, 257.7921, 258.5993, 259.7413, 260.5573, 
    260.7493, 259.3446, 256.2193, 250.8619, 261.405, 261.9633, 259.2309, 
    255.3995, 255.2062, 257.1832, 261.6096, 263.2114, 264.8473,
  271.3442, 272.7401, 272.9814, 273.1962, 273.0938, 272.8185, 272.4774, 
    272.2336, 270.3539, 270.5598, 270.4574, 270.1214, 269.3938, 268.0484, 
    266.6955, 266.5894, 267.4319, 268.4211, 269.2725, 270.0949,
  273.8025, 273.8303, 273.8063, 273.8644, 273.9276, 273.8366, 273.6484, 
    273.2454, 272.9586, 273.0345, 273.3212, 273.4842, 273.4084, 272.6012, 
    271.4807, 272.2727, 270.4018, 270.9551, 271.6209, 272.9094,
  274.6148, 274.755, 274.8434, 274.8144, 274.6641, 274.491, 274.4253, 
    274.6021, 274.9192, 275.3083, 275.5837, 275.7025, 275.7492, 275.6165, 
    275.3942, 275.2451, 275.1466, 275.0936, 274.9647, 274.9533,
  274.611, 274.8561, 275.3677, 275.662, 275.7505, 275.8566, 276.3, 276.6954, 
    276.9973, 277.0819, 276.8432, 276.5387, 276.5273, 276.7863, 276.9859, 
    277.116, 277.0339, 276.761, 276.2697, 275.9147,
  276.1761, 276.4301, 276.6082, 276.8242, 277.1375, 277.327, 277.4798, 
    277.7615, 277.639, 277.6137, 277.3725, 277.2133, 277.3636, 277.6706, 
    277.8651, 277.6213, 277.7666, 278.2769, 278.2883, 278.0395,
  278.618, 278.8985, 278.762, 278.6433, 278.7153, 278.8922, 279.1549, 
    279.0399, 278.9629, 278.7178, 278.5359, 278.6446, 278.9591, 279.1296, 
    279.453, 279.1322, 279.0109, 279.5832, 280.048, 280.1061,
  281.7926, 281.6776, 281.3542, 281.3466, 281.5677, 282.1134, 283.0482, 
    283.5245, 282.9447, 281.8191, 281.2683, 281.5968, 282.1059, 282.265, 
    282.596, 282.5606, 282.3244, 282.4621, 283.5637, 284.4037,
  284.8459, 284.4302, 284.4593, 285.0075, 286.2367, 288.3577, 290.6101, 
    291.555, 290.888, 288.9375, 287.481, 287.5303, 287.6996, 287.4355, 
    287.5303, 287.6301, 287.6402, 288.2326, 289.2205, 289.4744,
  287.5821, 287.6023, 287.956, 289.0032, 290.6101, 291.939, 293.3551, 
    295.0289, 296.037, 294.4592, 292.4127, 291.8114, 291.8961, 291.6813, 
    291.459, 291.6864, 292.0325, 291.891, 291.1179, 290.269,
  290.4181, 290.7806, 291.0939, 290.8716, 291.123, 288.4929, 289.3973, 
    291.9365, 293.11, 297.7424, 295.2942, 294.6449, 294.9316, 294.5779, 
    294.1472, 293.7025, 293.2819, 292.8675, 292.6047, 292.3546,
  292.8485, 293.1252, 292.4304, 291.1318, 290.989, 289.0197, 290.3852, 
    288.9919, 292.6805, 298.8932, 298.7694, 297.6754, 297.5238, 297.3811, 
    296.9668, 296.7836, 296.2328, 295.8374, 295.8905, 295.8829,
  294.0348, 293.3526, 292.3534, 291.6952, 290.9726, 291.6472, 292.0843, 
    288.412, 295.9637, 299.3202, 300.3422, 299.6878, 296.3099, 298.3892, 
    299.1105, 298.8035, 298.3854, 298.0557, 298.2729, 298.3702,
  294.8142, 293.9981, 293.8301, 295.3018, 292.7715, 292.0881, 292.8902, 
    294.0107, 296.3238, 298.6886, 301.5865, 301.5145, 292.6553, 294.4908, 
    299.7143, 299.7636, 299.5476, 299.3694, 299.559, 299.593,
  296.3958, 296.1052, 296.7507, 298.2628, 292.8827, 293.0166, 292.8384, 
    292.5706, 293.7354, 295.6959, 300.8816, 301.9553, 294.7649, 295.7187, 
    300.2083, 300.394, 300.4041, 300.418, 300.3485, 300.1287,
  251.2832, 250.8497, 250.4121, 250.0806, 249.6403, 249.2013, 248.7692, 
    248.3371, 247.8995, 247.3695, 246.9754, 246.5936, 246.209, 245.7524, 
    245.5241, 245.2292, 244.9615, 244.8596, 244.702, 244.6082,
  251.3172, 250.8348, 250.1635, 249.4052, 248.4988, 247.5584, 246.2403, 
    244.7794, 243.2615, 241.8958, 240.4105, 240.0518, 240.7516, 241.7966, 
    242.2546, 242.4869, 242.7098, 242.9435, 243.1378, 243.3267,
  252.6081, 251.3892, 250.6391, 249.9909, 249.2353, 248.5504, 248.208, 
    247.9389, 247.2268, 246.5922, 245.111, 243.7276, 243.6379, 243.3675, 
    243.5306, 243.5007, 243.7861, 244.2291, 244.5783, 246.084,
  247.4266, 243.0604, 239.5109, 236.0103, 232.9963, 236.827, 241.0329, 
    243.7942, 244.2182, 243.7399, 241.0506, 239.5068, 239.3356, 240.0721, 
    242.3225, 245.7782, 249.4378, 251.6922, 250.9856, 249.0111,
  260.4002, 254.584, 250.0479, 247.2758, 247.1806, 248.7774, 250.7043, 
    252.017, 252.5782, 252.5443, 251.2479, 250.3347, 250.5304, 250.7233, 
    250.7627, 251.5156, 253.2129, 256.0475, 257.3481, 257.0083,
  271.8083, 271.1098, 259.4109, 253.3868, 255.6535, 256.3751, 256.5137, 
    256.3615, 255.9932, 255.0311, 252.2738, 250.8647, 256.727, 255.0922, 
    250.5141, 247.0271, 253.149, 260.0849, 264.8995, 266.0736,
  273.0449, 272.4402, 271.9809, 271.7824, 271.9564, 270.9984, 270.7062, 
    270.3828, 270.1477, 272.114, 269.7794, 269.7278, 269.6177, 269.4981, 
    269.1516, 268.6936, 268.8214, 269.5416, 270.5064, 270.7538,
  275.6853, 275.0778, 274.4948, 274.2068, 274.0763, 274.0328, 274.0654, 
    273.8439, 273.5205, 273.3411, 273.3506, 273.3941, 273.4023, 272.8139, 
    271.8286, 272.3885, 269.774, 270.4453, 271.0391, 271.8993,
  275.2871, 274.9148, 274.696, 274.5845, 274.5397, 274.6172, 274.8264, 
    275.0629, 275.1308, 275.1335, 275.1036, 275.1403, 275.2844, 275.226, 
    274.8794, 274.4731, 274.2883, 274.4473, 274.7272, 275.5181,
  274.9052, 274.7408, 274.9229, 274.9827, 275.0425, 275.23, 275.6472, 
    275.9163, 276.1038, 276.2614, 276.3171, 276.3253, 276.5672, 276.858, 
    276.8023, 276.4612, 276.2248, 276.2886, 276.2424, 276.01,
  275.5045, 275.9747, 276.309, 276.449, 276.8906, 277.2942, 277.4315, 
    277.4899, 277.7807, 277.8799, 277.7821, 277.5157, 277.5864, 278.1395, 
    278.2386, 277.5578, 277.4451, 277.691, 277.865, 277.3812,
  278.3433, 278.6219, 278.5607, 278.3813, 278.5703, 278.7415, 278.6626, 
    278.7238, 278.8162, 278.6042, 278.4806, 278.6001, 278.7061, 278.7591, 
    278.7904, 278.5689, 278.3555, 278.5947, 279.2008, 278.9616,
  281.9186, 281.5422, 281.1291, 281.0122, 281.1318, 281.4172, 282.3834, 
    283.8782, 285.2221, 283.851, 282.5478, 282.204, 281.9526, 281.6074, 
    281.9037, 281.7963, 281.4892, 281.7053, 282.0803, 282.5097,
  284.6133, 284.0834, 284.0589, 284.2641, 285.252, 287.3733, 289.8329, 
    291.7843, 294.1815, 293.2954, 290.4458, 289.0461, 288.0745, 287.1477, 
    286.9466, 286.4587, 286.0144, 286.1285, 286.3215, 286.4397,
  287.4779, 287.3148, 287.2021, 287.675, 289.0679, 290.4879, 291.6634, 
    293.6732, 296.3843, 296.6859, 294.5416, 293.3349, 292.5766, 291.4351, 
    290.6035, 289.8574, 289.341, 289.4239, 289.394, 289.3967,
  290.5355, 290.2094, 290.0191, 290.1917, 290.0341, 285.5184, 285.1447, 
    284.6582, 293.7031, 298.583, 296.2783, 295.876, 296.3802, 294.5973, 
    293.8173, 293.5251, 293.021, 292.7111, 292.7166, 292.7763,
  292.3727, 292.0453, 291.5248, 291.2843, 290.0775, 282.4825, 284.5277, 
    287.6994, 293.627, 299.5587, 298.9091, 297.9226, 297.8125, 297.6032, 
    297.2526, 297.0461, 296.3204, 295.7293, 295.7945, 295.9603,
  293.4694, 293.0046, 292.2559, 291.4894, 285.9424, 285.483, 290.2189, 
    291.9053, 293.9083, 297.9769, 301.2601, 300.3672, 296.7403, 298.6374, 
    299.1809, 298.5721, 298.0381, 297.8573, 298.2596, 298.3982,
  294.8867, 294.1774, 294.0796, 295.2795, 287.2034, 290.3548, 293.7955, 
    293.9586, 293.7004, 295.0811, 302.3146, 301.7615, 294.3078, 294.5484, 
    299.6783, 299.8468, 299.5927, 299.4242, 299.5193, 299.3888,
  296.5433, 295.9684, 296.5147, 298.2066, 290.6143, 291.8414, 294.1815, 
    293.5577, 292.9095, 295.7252, 301.983, 301.6935, 294.8949, 295.1245, 
    300.0764, 300.4923, 300.283, 300.1376, 299.9881, 299.8101 ;
}
