netcdf tnhus_cfSites_exAA04_amip_r3i1p1_1998_slice {
dimensions:
	site = 120 ;
	mlev = 62 ;
	nhym = 62 ;
	nhyi = 63 ;
	time = UNLIMITED ; // (10 currently)
variables:
	double site(site) ;
		site:standard_name = "latitude" ;
		site:long_name = "site index" ;
		site:units = "degrees_north" ;
		site:axis = "Y" ;
	double mlev(mlev) ;
		mlev:standard_name = "hybrid_sigma_pressure" ;
		mlev:long_name = "hybrid level at layer midpoints" ;
		mlev:formula = "hyam hybm (mlev=hyam+hybm*aps)" ;
		mlev:formula_terms = "ap: hyam b: hybm ps: aps" ;
		mlev:units = "level" ;
		mlev:positive = "down" ;
	double hyai(nhyi) ;
		hyai:long_name = "hybrid A coefficient at layer interfaces" ;
		hyai:units = "Pa" ;
	double hybi(nhyi) ;
		hybi:long_name = "hybrid B coefficient at layer interfaces" ;
		hybi:units = "1" ;
	double hyam(nhym) ;
		hyam:long_name = "hybrid A coefficient at layer midpoints" ;
		hyam:units = "Pa" ;
	double hybm(nhym) ;
		hybm:long_name = "hybrid B coefficient at layer midpoints" ;
		hybm:units = "1" ;
	double time(time) ;
		time:standard_name = "time" ;
		time:units = "hours since 1998-1-1 03:00:00" ;
		time:calendar = "proleptic_gregorian" ;
		time:axis = "T" ;
	float tnhus(time, mlev, site) ;
		tnhus:long_name = "Tendency of Air Temperature" ;
		tnhus:units = "K s**-1" ;
		tnhus:table = 128 ;
		tnhus:grid_type = "gaussian" ;

// global attributes:
		:CDI = "Climate Data Interface version ?? (http://mpimet.mpg.de/cdi)" ;
		:Conventions = "CF-1.0" ;
		:history = "reset by cdo to create anonymous sample file" ;
		:source = "201707_compliance_checker_evaluation/work/p1.py" ;
		:institution = "CEDA" ;
		:product = "output" ;
		:physics_version = 1 ;
		:references = "Model described by Hazeleger et al. (Bull. Amer. Meteor. Soc., 2010, 91, 1357-1363). Also see http://ecearth.knmi.nl" ;
		:freqency = "subhr" ;
		:title = "Dummy file with known metadata errors" ;
		:contact = "none" ;
		:realization = 3 ;
		:project_id = "CMIP5" ;
		:institute_id = "CEDA" ;
		:initialization_method = 1 ;
		:parent_experiment_id = "N/A" ;
		:creation_date = "2013-02-20T20:10:51Z2013-02-24T12:00" ;
		:parent_experiment = "piControl" ;
		:branch_time = 0 ;
		:forcing = "Nat,Ant" ;
		:modeling_realm = "atmos" ;
		:table_id = "Table cfSites (01 February 2012) 69520b77c6b6f66ea514a9e1ed36acfb" ;
		:experiment_id = "amip" ;
		:parent_experiment_rip = "N/A" ;
		:tracking_id = "04190a74-1606-49d7-9d2d-89bc32058df6" ;
		:model_id = "exAA04" ;
		:frequency = "subhr" ;
		:comment = "this is a sample file with known metadata errors" ;
		:CDO = "Climate Data Operators version 1.7.0 (http://mpimet.mpg.de/cdo)" ;
data:

 site = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 
    20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 37, 
    38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 55, 
    56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 72, 73, 
    74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 90, 91, 
    92, 93, 94, 95, 96, 97, 98, 99, 100, 101, 102, 103, 104, 105, 106, 107, 
    108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 120 ;

 mlev = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 
    20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 37, 
    38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 55, 
    56, 57, 58, 59, 60, 61, 62 ;

 hyai = 0, 988.8359375, 1977.67626953125, 2966.5166015625, 3955.35693359375, 
    4944.19921875, 5933.0390625, 6921.87109375, 7909.44140625, 8890.70703125, 
    9860.52734375, 10807.78125, 11722.75, 12595.0078125, 13419.46484375, 
    14192.01171875, 14922.6875, 15638.0546875, 16329.5625, 16990.625, 
    17613.28125, 18191.03125, 18716.96875, 19184.546875, 19587.515625, 
    19919.796875, 20175.39453125, 20348.91796875, 20434.15625, 20426.21875, 
    20319.01171875, 20107.03125, 19785.359375, 19348.77734375, 
    18798.82421875, 18141.296875, 17385.59375, 16544.5859375, 15633.56640625, 
    14665.64453125, 13653.21875, 12608.3828125, 11543.16796875, 10471.3125, 
    9405.22265625, 8356.25390625, 7335.1640625, 6353.921875, 5422.80078125, 
    4550.21484375, 3743.46435546875, 3010.14697265625, 2356.20263671875, 
    1784.8544921875, 1297.65625, 895.193603515625, 576.314208984375, 
    336.7724609375, 162.043426513672, 54.2083435058594, 6.57562828063965, 
    0.00316000008024275, 0 ;

 hybi = 0, 0, 0, 0, 0, 0, 0, 7.59000045036373e-08, 1.25998003568384e-05, 
    8.73560929903761e-05, 0.00027506984770298, 0.000685490202158689, 
    0.00141457631252706, 0.0025651603937149, 0.00418749824166298, 
    0.00632216781377792, 0.00903499126434326, 0.0125082619488239, 
    0.0168595798313618, 0.0221886448562145, 0.0286103487014771, 
    0.0362269096076488, 0.0451461337506771, 0.055474229156971, 
    0.0673161745071411, 0.0807772874832153, 0.0959640741348267, 
    0.112978994846344, 0.131934821605682, 0.152933537960052, 
    0.176091074943542, 0.201520144939423, 0.229314863681793, 
    0.259554445743561, 0.29199343919754, 0.326329410076141, 0.3622025847435, 
    0.399204790592194, 0.436906337738037, 0.475016415119171, 
    0.513279736042023, 0.551458477973938, 0.589317142963409, 
    0.626558899879456, 0.662933588027954, 0.69822359085083, 
    0.732223808765411, 0.764679491519928, 0.795384764671326, 
    0.824185431003571, 0.850950419902802, 0.875518381595612, 
    0.897767245769501, 0.917650938034058, 0.935157060623169, 
    0.950273811817169, 0.963007092475891, 0.973466038703918, 
    0.982238113880157, 0.98915296792984, 0.994204163551331, 0.99763011932373, 1 ;

 hyam = 494.41796875, 1483.25610351562, 2472.09643554688, 3460.93676757812, 
    4449.77807617188, 5438.619140625, 6427.455078125, 7415.65625, 
    8400.07421875, 9375.6171875, 10334.154296875, 11265.265625, 
    12158.87890625, 13007.236328125, 13805.73828125, 14557.349609375, 
    15280.37109375, 15983.80859375, 16660.09375, 17301.953125, 17902.15625, 
    18454, 18950.7578125, 19386.03125, 19753.65625, 20047.595703125, 
    20262.15625, 20391.537109375, 20430.1875, 20372.615234375, 
    20213.021484375, 19946.1953125, 19567.068359375, 19073.80078125, 
    18470.060546875, 17763.4453125, 16965.08984375, 16089.076171875, 
    15149.60546875, 14159.431640625, 13130.80078125, 12075.775390625, 
    11007.240234375, 9938.267578125, 8880.73828125, 7845.708984375, 
    6844.54296875, 5888.361328125, 4986.5078125, 4146.83959960938, 
    3376.8056640625, 2683.1748046875, 2070.52856445312, 1541.25537109375, 
    1096.42492675781, 735.75390625, 456.543334960938, 249.407943725586, 
    108.125885009766, 30.3919858932495, 3.28939414035995, 0.00158000004012138 ;

 hybm = 0, 0, 0, 0, 0, 0, 3.79500022518187e-08, 6.33785018067101e-06, 
    4.99779466736072e-05, 0.000181212970346678, 0.000480280024930835, 
    0.00105003325734288, 0.00198986835312098, 0.00337632931768894, 
    0.00525483302772045, 0.00767857953906059, 0.0107716266065836, 
    0.0146839208900928, 0.0195241123437881, 0.0253994967788458, 
    0.032418629154563, 0.040686521679163, 0.050310181453824, 
    0.061395201832056, 0.0740467309951782, 0.088370680809021, 
    0.104471534490585, 0.122456908226013, 0.142434179782867, 
    0.164512306451797, 0.188805609941483, 0.215417504310608, 
    0.244434654712677, 0.275773942470551, 0.309161424636841, 
    0.344265997409821, 0.380703687667847, 0.418055564165115, 
    0.455961376428604, 0.494148075580597, 0.53236910700798, 
    0.570387810468674, 0.607938021421432, 0.644746243953705, 
    0.680578589439392, 0.715223699808121, 0.74845165014267, 
    0.780032128095627, 0.809785097837448, 0.837567925453186, 
    0.863234400749207, 0.886642813682556, 0.907709091901779, 
    0.926403999328613, 0.942715436220169, 0.95664045214653, 
    0.968236565589905, 0.977852076292038, 0.985695540904999, 
    0.991678565740585, 0.995917141437531, 0.998815059661865 ;

 time = 0, 3, 6, 9, 12, 15, 18, 21, 24, 27 ;

 tnhus =
  6.179532e-13, 2.689177e-13, 5.555486e-14, -8.39057e-14, -2.302788e-13, 
    -2.748213e-13, -1.390936e-13, 1.334925e-13, 5.842923e-13, 5.605742e-13, 
    -4.8459e-14, -3.448012e-13, -4.504902e-14, 1.476382e-13, 1.939659e-14, 
    6.692602e-13, 4.972176e-14, -5.505814e-12, -5.129654e-14, -6.606461e-14, 
    -4.506272e-13, -3.13143e-12, -1.076993e-12, 3.789546e-13, -2.257472e-13, 
    -3.815103e-13, -6.823792e-14, -7.954256e-14, -1.652043e-13, 1.83527e-14, 
    -4.496357e-14, -7.778118e-14, -5.043799e-14, -4.766506e-14, 
    -1.031724e-13, -6.863427e-14, 2.713804e-14, 4.776018e-13, 1.70832e-13, 
    1.204367e-13, 7.058703e-13, 1.246433e-12, -1.694364e-14, -7.86775e-15, 
    1.651737e-13, 3.776412e-15, 2.044235e-14, 4.558969e-14, 2.161964e-12, 
    1.388185e-12, 4.543156e-13, -7.524094e-13, -7.777207e-13, -4.970306e-13, 
    3.128476e-13, -7.617961e-13, -9.595758e-15, 9.906673e-13, -1.440525e-13, 
    -1.112811e-12, 9.013978e-13, 1.304552e-12, 4.145555e-13, -7.41606e-13, 
    -3.042281e-12, -1.98695e-13, 2.298021e-13, 8.004685e-14, 6.152449e-14, 
    1.653416e-13, 4.237815e-13, 9.689813e-14, -2.291759e-13, 2.333255e-14, 
    4.847824e-14, -7.508713e-13, 6.343315e-13, -1.941539e-13, -3.087414e-12, 
    -1.422239e-12, 3.109544e-13, -1.776989e-12, 5.778931e-13, -3.223701e-13, 
    -3.203613e-13, 4.694089e-14, 3.675027e-13, -3.309904e-13, 4.171754e-13, 
    6.231963e-13, -2.386988e-14, 9.465005e-13, 4.298002e-14, 1.624702e-13, 
    -3.618918e-15, 2.708928e-14, 2.128039e-13, -2.542991e-13, -3.701102e-13, 
    -1.586456e-13, 3.582297e-13, 4.073472e-13, -5.549118e-14, 4.496655e-13, 
    5.041823e-14, -9.901016e-15, -2.079522e-13, -7.21489e-14, -5.696803e-14, 
    -3.975893e-14, 5.590535e-14, 1.779109e-14, 4.770291e-13, 4.926293e-13, 
    9.195382e-13, -4.453515e-12, 8.839513e-13, 2.779061e-13, 4.875848e-13, 
    -1.387504e-12,
  -1.124503e-13, -1.178959e-13, -8.138547e-14, 3.706619e-14, 1.142157e-13, 
    1.557459e-13, 3.078653e-13, 4.395413e-13, 3.808106e-13, 2.74425e-13, 
    7.983114e-14, 8.773642e-14, -1.411983e-13, 3.817104e-13, 6.75268e-13, 
    2.114166e-14, -1.123161e-13, -1.177012e-13, 1.866079e-13, 2.891644e-13, 
    1.639765e-13, 1.953465e-12, 2.990961e-12, 6.86974e-14, 5.110084e-14, 
    1.937668e-13, 4.613627e-14, -2.073943e-13, -1.223476e-13, -1.366971e-13, 
    -9.359145e-14, -2.106821e-13, -8.085762e-14, 2.177964e-15, -5.298716e-14, 
    3.451413e-14, -1.464371e-12, 6.159601e-13, -2.236216e-13, 1.787864e-12, 
    3.428273e-13, -2.595852e-13, 2.384555e-13, 1.543273e-13, 2.184656e-13, 
    8.266356e-13, -6.339961e-13, -1.294833e-13, 1.760174e-13, -7.304887e-13, 
    2.483879e-13, -4.53847e-13, 6.978436e-14, -9.515544e-12, 5.381428e-13, 
    -1.056642e-12, 1.271426e-13, -5.888814e-13, 5.455454e-13, 1.334161e-12, 
    3.016671e-13, -1.900367e-13, -3.133785e-13, -8.010164e-14, -7.696552e-14, 
    -2.108554e-14, 3.755239e-13, 4.817476e-13, 1.067039e-13, 4.946038e-14, 
    6.08534e-13, 1.573439e-13, 4.323154e-13, -9.773674e-14, -2.33019e-14, 
    -2.119809e-13, -3.682833e-13, -1.524393e-13, 7.082476e-12, -3.255551e-12, 
    -1.805543e-13, 3.915424e-13, 1.588109e-12, 3.012839e-13, -2.628599e-13, 
    -2.864503e-13, 6.809495e-13, -3.891027e-13, 1.542173e-12, 3.687775e-13, 
    -2.546319e-13, -1.105203e-12, -4.764355e-14, 3.727903e-14, -4.990433e-14, 
    6.326385e-13, -1.847066e-13, 2.633324e-13, 8.959716e-13, -7.75091e-13, 
    -8.604193e-13, 1.530864e-13, -5.914942e-13, 6.766294e-14, -6.710319e-13, 
    2.694354e-13, 7.430134e-14, -1.016759e-12, -2.326383e-13, -1.639447e-13, 
    -3.221974e-14, 2.383223e-13, 2.089027e-13, 5.510831e-13, 1.695239e-13, 
    -9.291433e-13, -1.799186e-13, 2.518166e-12, -6.095303e-14, -9.972478e-14,
  -2.149947e-13, -2.355338e-13, -9.003909e-14, 1.497413e-14, -1.484923e-15, 
    -8.223977e-14, -8.504308e-14, -6.175616e-15, -2.920858e-13, 
    -4.425627e-14, 4.744816e-14, 3.777534e-14, -1.321443e-13, -6.926404e-14, 
    -1.733474e-13, -1.592129e-13, -2.634906e-13, -3.204173e-13, 
    -5.907826e-13, -1.085451e-12, -2.97512e-13, -8.031076e-13, -9.871548e-13, 
    -3.463618e-13, -9.663104e-13, -5.805495e-13, -1.283418e-13, 
    -3.935463e-13, -4.638651e-13, -3.465839e-13, -2.47441e-13, -1.729172e-13, 
    -7.659151e-14, 5.040413e-14, -4.249379e-14, -1.078165e-13, -9.452439e-13, 
    -1.851297e-14, 1.167955e-13, 3.810452e-13, -6.138784e-13, 4.562323e-13, 
    -4.163579e-13, -7.675913e-14, 5.073719e-14, 7.909506e-13, -1.646093e-12, 
    -5.721812e-13, -1.750061e-12, -9.430737e-14, -1.571313e-14, 
    -4.430345e-13, -2.666437e-13, -3.326095e-12, 2.004646e-14, -1.61382e-12, 
    -8.441303e-13, -5.89942e-13, 1.014079e-12, -8.613249e-14, -2.513961e-13, 
    8.769097e-13, -5.121459e-13, -2.55404e-13, -6.019046e-13, 2.975536e-13, 
    -1.570688e-13, -4.755918e-14, -8.439083e-14, -2.042533e-13, 2.319228e-12, 
    2.7639e-13, -5.241363e-13, 6.620815e-13, -2.34314e-13, -1.43989e-12, 
    -1.771812e-13, 8.424025e-13, -2.56225e-12, -1.68629e-13, 6.812745e-13, 
    5.95584e-13, -4.387324e-13, -3.685108e-13, 2.733924e-14, -5.922624e-13, 
    -1.323552e-12, 9.925394e-14, 6.219227e-13, -1.031536e-13, -6.136758e-14, 
    -1.362577e-13, 4.2958e-13, -4.518594e-13, 1.074141e-14, 7.588235e-14, 
    -4.30922e-13, 2.665923e-14, 3.901324e-13, -3.348516e-13, -2.139955e-14, 
    4.718066e-13, -3.312654e-13, -3.904689e-14, -3.269884e-13, 7.907563e-13, 
    1.064857e-12, 1.595987e-12, 1.761521e-12, 1.111694e-12, 1.089545e-12, 
    6.882411e-13, 7.529394e-13, 4.978934e-13, -5.783707e-13, -9.626438e-13, 
    5.268438e-12, 6.160263e-12, -9.851495e-13, 4.991979e-13,
  -2.660511e-13, -3.26475e-13, -2.664674e-13, -1.671996e-13, -9.486856e-14, 
    -5.707934e-14, -1.242617e-13, -1.669498e-14, 5.094536e-14, 4.296563e-13, 
    3.574918e-13, 2.287337e-13, 3.2363e-13, 1.445649e-13, 3.812783e-13, 
    -3.243364e-13, -1.296796e-13, -3.884948e-13, -3.854451e-13, 
    -5.417611e-13, -2.160772e-13, -1.958295e-13, -3.698986e-13, 
    -7.444462e-13, -2.706307e-13, -2.595146e-13, -2.326611e-13, 8.476553e-14, 
    1.092043e-13, 2.40169e-13, -8.149037e-14, 2.042949e-13, 4.000827e-13, 
    -1.077194e-13, 3.219647e-15, -2.385453e-13, -8.613804e-14, -7.297253e-13, 
    -1.424e-13, 1.115098e-12, 1.588979e-13, -5.226791e-13, -6.24896e-13, 
    -2.307551e-13, 2.412931e-13, 1.681308e-12, 1.29434e-12, 1.501559e-12, 
    -1.560696e-14, 1.538651e-11, 1.782104e-12, -1.614014e-12, -7.855564e-13, 
    -2.370881e-14, 2.763858e-13, -4.061196e-13, -1.696213e-12, -1.829842e-12, 
    5.743475e-13, 1.121197e-12, 6.159934e-13, 1.271205e-13, 6.641632e-13, 
    -2.121359e-13, -2.028599e-13, -1.244893e-12, -8.315848e-13, 
    -5.044853e-13, -2.161465e-13, -2.365746e-13, 8.782142e-13, -6.415563e-13, 
    -1.825484e-13, -9.214851e-15, -3.222922e-13, -1.281197e-12, 
    -1.092628e-12, 2.068297e-12, -2.922572e-11, 8.651413e-14, 9.211382e-13, 
    1.728102e-12, 2.856743e-14, 2.400163e-13, -1.063039e-14, -2.863682e-13, 
    -1.060541e-13, 4.277273e-13, 1.304125e-12, -1.746339e-12, -1.441625e-13, 
    -1.287492e-12, 1.089875e-12, 6.909112e-13, 2.355477e-13, -4.002354e-14, 
    -1.701139e-14, -2.040035e-13, -6.299544e-13, -1.094891e-12, 1.054545e-12, 
    7.134397e-14, 6.546222e-13, -2.723707e-13, 1.908335e-13, 4.815731e-13, 
    7.541329e-13, 9.100637e-13, 5.416778e-13, 5.845324e-14, -3.302913e-14, 
    2.036843e-13, 5.991041e-14, 7.571721e-14, 2.302186e-13, 1.450717e-12, 
    1.566211e-11, -1.201085e-11, 3.220132e-13, 8.050227e-13,
  -2.855494e-13, -4.282408e-13, -4.929945e-13, -5.19057e-13, -4.239109e-13, 
    -3.350098e-13, 9.88376e-14, -7.244205e-15, -2.813305e-13, 1.417144e-12, 
    -1.057765e-13, 6.095124e-14, -1.323941e-13, -1.523781e-13, -2.050304e-13, 
    -3.414852e-13, -2.149197e-13, -6.041417e-13, -8.859406e-13, 
    -6.440404e-13, -7.589762e-13, -1.332101e-12, -4.058698e-13, -1.75443e-13, 
    -4.512779e-13, -1.544598e-13, 1.117439e-13, -6.944445e-14, -2.181588e-13, 
    2.012279e-14, -2.046086e-12, -5.58914e-13, 5.489498e-13, 9.835743e-13, 
    -4.103384e-13, -5.832834e-13, -1.850853e-13, 1.440088e-12, -4.610201e-14, 
    -1.6385e-12, 1.380285e-12, -1.469658e-13, -7.73312e-13, -4.590061e-13, 
    2.232492e-12, 1.300182e-12, 5.704742e-13, 2.415831e-12, 8.830381e-13, 
    2.446529e-11, 1.277908e-12, -2.390588e-12, 3.770284e-12, 5.111412e-13, 
    1.925946e-13, -5.462436e-13, -3.004763e-12, 1.264913e-12, 5.69303e-13, 
    2.88242e-12, -1.043082e-12, -3.438083e-13, -5.840051e-13, -2.684852e-13, 
    -4.669154e-13, -3.826106e-13, 2.670364e-13, 3.198553e-13, 7.912837e-13, 
    1.081774e-12, -1.070533e-13, -4.177214e-13, -1.179001e-12, -1.041389e-13, 
    -8.213375e-13, -9.82936e-13, 1.170203e-12, -4.559339e-13, 2.344179e-12, 
    -3.014256e-14, 1.103825e-12, 1.452816e-12, 6.902812e-14, -4.397593e-13, 
    2.009504e-14, 2.088607e-13, -3.869127e-14, -4.624912e-13, -1.233489e-12, 
    2.939538e-12, -4.751755e-13, 9.22229e-13, 3.468406e-13, 1.61752e-12, 
    4.951595e-14, 5.65521e-12, 4.757833e-12, -3.744505e-13, -1.000205e-11, 
    8.879564e-13, 1.629946e-12, 4.259353e-13, 1.121105e-12, -1.439734e-13, 
    -3.077538e-13, 2.810252e-13, 2.433054e-13, -3.559375e-13, -9.033885e-13, 
    -1.031425e-12, -8.233136e-13, -8.012757e-13, -4.757861e-13, 
    -4.123646e-13, -5.305201e-13, 6.277367e-13, 3.230537e-12, -2.676089e-11, 
    -5.958289e-13, -3.104184e-13,
  -2.187833e-13, -4.105188e-13, -5.205697e-13, -3.747419e-13, -4.821282e-13, 
    -5.244416e-14, 2.757378e-13, 6.23876e-13, 4.126283e-13, -4.938411e-13, 
    2.041284e-13, -4.463235e-13, -5.902917e-13, -1.314324e-12, 1.380493e-12, 
    -3.170353e-13, -1.424e-12, -1.713366e-12, -7.801156e-13, -5.491302e-13, 
    -3.293338e-13, 1.384864e-13, -1.790804e-12, -2.467568e-12, -6.185746e-13, 
    -1.530456e-12, -1.428066e-12, -1.215514e-12, -1.183678e-12, 
    -8.928552e-13, 4.69666e-13, 7.950446e-13, -1.214723e-13, -9.395401e-13, 
    -5.825479e-13, 5.326434e-13, -5.393463e-14, 6.839928e-12, -3.265027e-13, 
    5.221132e-12, -2.456785e-13, -1.419961e-12, -1.361231e-12, -1.223794e-12, 
    -2.344611e-12, 3.205672e-12, 8.721218e-13, -5.126524e-13, 1.938255e-13, 
    1.428835e-11, -4.424308e-13, 7.320394e-13, -5.132283e-13, 7.609561e-12, 
    4.676696e-13, 6.790263e-13, 1.263226e-12, 6.429079e-13, 4.331951e-13, 
    5.761974e-12, -1.003295e-12, 7.840534e-13, -1.404085e-12, -7.678719e-13, 
    -1.551978e-12, 4.779371e-13, -4.349437e-13, -1.208519e-12, -1.007801e-11, 
    -8.329032e-13, -8.012063e-13, 9.37958e-13, -1.472475e-12, -4.723028e-13, 
    -4.703987e-13, -1.290815e-12, 8.216344e-14, -3.455639e-13, -8.104669e-12, 
    -2.597991e-12, 1.690342e-12, 1.753583e-13, 1.475764e-13, -4.005823e-13, 
    7.320533e-14, 5.24368e-12, 2.85634e-12, -5.116602e-13, -5.34634e-13, 
    2.77775e-12, -1.116482e-12, -3.310324e-13, -9.747134e-13, 8.332252e-13, 
    7.846918e-13, 2.726436e-12, 8.430451e-13, 1.274397e-13, -5.495174e-12, 
    -2.638528e-13, 3.328379e-12, 2.032673e-12, 1.533079e-13, -7.682396e-13, 
    -4.804074e-13, -8.718443e-13, -1.167108e-12, -1.474834e-12, 
    -1.460818e-12, -1.189257e-12, -1.05653e-12, -1.563596e-12, -6.124407e-13, 
    -2.974704e-13, 1.078984e-12, 4.929834e-13, -1.351844e-11, 2.795948e-12, 
    5.093755e-13, 6.973588e-14,
  -2.305378e-13, 3.538281e-13, 4.267697e-13, 6.243339e-13, 1.981804e-12, 
    -4.536926e-13, 1.121603e-12, -2.441936e-13, -8.48932e-13, 4.04532e-12, 
    3.48771e-12, 2.594425e-12, -2.865264e-12, -7.141066e-12, 4.657386e-13, 
    -1.892891e-12, -3.700884e-12, 1.717265e-12, -4.130613e-12, -3.511247e-12, 
    -5.919709e-13, 1.604272e-13, -1.025957e-12, -2.308209e-12, -3.000766e-12, 
    -5.237699e-12, -6.919298e-12, -9.255818e-12, -1.070849e-11, 
    -8.814838e-12, -2.669975e-12, 6.305345e-12, 5.314416e-12, -9.204859e-13, 
    1.976752e-12, -4.166167e-12, 1.861455e-13, 4.845409e-12, -8.926193e-14, 
    1.424472e-13, 2.092371e-12, 2.712719e-12, -4.250642e-12, -1.897493e-12, 
    3.601008e-13, 4.721001e-12, 3.854306e-12, 1.758732e-13, 2.588607e-12, 
    -1.274104e-11, 2.164588e-13, 1.790568e-12, 3.333833e-13, 7.17626e-12, 
    9.733825e-13, 3.300971e-13, 1.282086e-12, 1.647488e-12, 2.609096e-12, 
    5.619498e-12, 5.400791e-12, 8.030243e-13, -1.495859e-12, -1.965661e-12, 
    -3.50765e-12, 1.234013e-12, -1.82182e-12, 9.286627e-12, 8.399947e-12, 
    9.711676e-12, -3.417933e-12, 1.29054e-11, -3.31063e-12, 6.332712e-13, 
    4.72028e-13, -1.931788e-14, -8.442552e-14, 1.698391e-12, -8.404605e-12, 
    2.274181e-12, 4.225592e-12, 8.127272e-12, 1.951495e-13, -7.426948e-12, 
    -1.766476e-12, 5.828282e-12, 1.411232e-11, -8.392176e-13, 4.169196e-12, 
    -7.786272e-13, 1.03384e-12, -6.38134e-13, 3.47361e-14, -3.996331e-12, 
    4.542144e-12, -5.781253e-12, -2.774592e-12, -1.495137e-12, 1.068312e-11, 
    1.473843e-12, 1.017131e-12, 1.957202e-12, -2.08282e-12, -3.163124e-11, 
    -2.610689e-13, -2.225942e-12, -3.543998e-12, -1.52367e-12, -1.860567e-12, 
    -3.6392e-12, -3.98781e-12, 7.421286e-13, -4.060086e-13, 2.229883e-13, 
    -1.084133e-13, 4.894196e-13, -1.104533e-13, -3.039635e-12, 2.279496e-13, 
    1.938893e-12,
  -4.855838e-13, -5.499406e-12, -1.439943e-11, -1.802014e-11, -1.377529e-11, 
    -1.079634e-11, -4.226314e-12, -4.082151e-12, -7.338158e-12, 
    -8.317902e-12, -1.011211e-11, 1.007586e-11, 1.690037e-12, 1.824652e-12, 
    -8.528206e-12, -1.016892e-12, 3.893375e-12, -2.703324e-12, -7.772092e-12, 
    3.043676e-13, 1.431077e-12, 2.797762e-14, 3.3476e-13, -4.271306e-13, 
    -1.979222e-12, -2.744194e-13, -1.059614e-11, -4.650558e-12, 
    -5.904499e-12, -1.160264e-11, 3.868267e-12, 6.630502e-12, 7.68452e-12, 
    1.155992e-12, 3.839568e-12, 3.437667e-12, -9.141937e-13, 9.739119e-13, 
    7.861795e-12, 6.898204e-13, -1.929286e-11, 3.138989e-12, 1.214959e-12, 
    -1.07155e-12, -2.398776e-12, 2.373463e-12, 6.053005e-12, 6.508682e-14, 
    1.404232e-12, -2.952208e-12, 4.867516e-12, 1.703498e-12, 9.02009e-13, 
    3.878009e-14, 7.544035e-13, 1.637718e-13, 8.245182e-12, 6.769721e-12, 
    3.438258e-12, 3.0888e-12, 1.937422e-12, 2.366107e-12, -3.190337e-12, 
    4.559092e-12, 4.256995e-12, -7.340212e-12, 1.515205e-11, 1.823869e-11, 
    2.195691e-11, -4.711703e-12, 4.751199e-13, -9.591328e-12, -4.419909e-12, 
    -1.134481e-12, 2.14733e-12, -5.022094e-13, -2.096379e-13, 8.180887e-13, 
    2.910183e-12, 1.052303e-11, 6.011358e-12, 9.853281e-12, 1.866757e-12, 
    -1.946682e-11, -3.452794e-13, 1.524364e-12, 1.310513e-11, 4.832745e-12, 
    -4.721189e-13, 6.976641e-13, 8.049117e-14, 1.440237e-13, 2.790823e-14, 
    2.935413e-12, -1.914802e-12, -1.164602e-11, 1.428774e-12, -1.133849e-11, 
    6.189271e-12, 3.903833e-12, -8.334805e-12, 7.97782e-13, -5.725854e-13, 
    -3.037149e-11, -1.066508e-12, -1.612349e-12, -3.425621e-12, 
    -3.457151e-12, -3.261641e-12, -4.459016e-12, -6.599443e-13, -5.93614e-12, 
    -6.008943e-12, -4.808931e-12, -1.884298e-12, 1.151884e-12, 1.590884e-12, 
    -2.58504e-12, 9.307659e-14, 2.996797e-12,
  -8.18709e-12, -2.420167e-11, -1.890532e-11, -1.357806e-11, -1.627137e-11, 
    -1.460423e-11, -9.127865e-12, -2.318287e-11, 2.70039e-11, 2.314005e-11, 
    -1.062095e-12, 2.600142e-13, -9.714451e-14, -3.158696e-12, -5.164591e-12, 
    5.813014e-12, 2.661538e-12, -9.102857e-12, -1.030592e-12, -9.449108e-13, 
    1.454142e-12, -1.864814e-12, -3.756273e-12, -5.641848e-12, -4.532569e-12, 
    -1.249001e-15, -6.102896e-13, -1.14303e-11, 3.012363e-11, 6.083023e-12, 
    4.534983e-12, -5.76908e-12, -4.453105e-13, 2.890743e-12, 2.218675e-11, 
    -2.688191e-11, -2.639744e-12, 2.619693e-12, -1.363432e-11, 3.71691e-12, 
    2.999451e-12, 1.859901e-12, 3.568257e-13, -2.475232e-12, -5.543455e-12, 
    3.426981e-12, 5.29353e-12, -7.192233e-13, 1.283129e-12, 2.159959e-11, 
    6.772735e-12, -2.011447e-13, 2.004349e-12, 1.022665e-12, 4.496063e-13, 
    9.680312e-13, 4.546363e-14, 8.867548e-12, 1.966419e-12, 1.487578e-11, 
    -4.317657e-12, 4.347439e-12, -1.448813e-12, 5.534112e-12, 1.157602e-12, 
    2.575523e-12, 2.949938e-11, 1.166087e-11, 3.893996e-12, -3.120293e-11, 
    4.444306e-12, 3.501643e-13, 4.480583e-13, -1.628142e-11, -1.984379e-12, 
    -5.701134e-12, -5.992429e-13, 1.852823e-13, 1.602922e-11, 3.078093e-13, 
    6.62953e-12, -3.515357e-12, 1.698044e-12, -1.905218e-11, -6.57091e-12, 
    -4.188705e-12, -1.22754e-11, -1.20853e-11, -2.918624e-12, 2.874284e-12, 
    4.657164e-12, -3.822687e-12, -3.637229e-13, 6.551457e-12, -1.41348e-12, 
    -1.106681e-11, -2.026385e-12, 1.086677e-10, -3.969325e-13, 1.755973e-12, 
    -8.118645e-12, 6.162557e-12, 6.965244e-13, -1.399888e-11, 3.305106e-12, 
    4.55358e-13, -1.947248e-12, -8.098494e-12, -1.064057e-11, -3.518019e-13, 
    -3.581385e-12, -1.024442e-11, -1.594355e-11, -1.43684e-11, 7.939538e-12, 
    9.875767e-13, 1.808866e-13, -2.110141e-12, -9.074547e-13, 3.09644e-12,
  -1.347711e-11, -1.648581e-11, -1.02256e-11, -3.052891e-12, -8.437473e-12, 
    -4.812928e-12, -8.625989e-12, 8.263268e-11, 1.54548e-10, 6.667922e-11, 
    1.51521e-11, -3.47633e-12, -6.919687e-12, -1.79412e-11, -1.373368e-11, 
    5.574186e-12, -6.691314e-14, -1.304079e-11, -6.840445e-12, -9.665602e-13, 
    -1.602163e-12, -1.661438e-11, -1.983969e-12, -2.10667e-11, 5.716538e-13, 
    1.853284e-11, -1.949252e-11, -4.441447e-12, 1.388845e-11, -2.917599e-11, 
    3.816725e-11, -1.654488e-11, 2.390999e-11, -5.010437e-12, 6.939327e-11, 
    -1.334751e-10, -9.003554e-12, 3.422984e-12, -5.29834e-11, 4.059708e-12, 
    1.518825e-11, -1.82343e-12, -2.284478e-12, -1.747422e-12, 2.63578e-12, 
    5.514367e-12, 2.069345e-12, -1.051853e-12, 1.355938e-12, 1.139181e-11, 
    1.152647e-12, -5.219047e-12, 2.208123e-12, 1.20759e-12, 5.99501e-13, 
    1.000533e-12, -3.824763e-11, 8.494904e-12, -2.915313e-12, 2.873109e-11, 
    -1.516887e-11, 1.09901e-11, 7.805534e-12, 4.348766e-12, -2.539924e-12, 
    -1.150898e-10, -4.846457e-12, 3.295808e-12, 5.02306e-11, -1.482492e-11, 
    -6.726841e-13, 2.044032e-12, 1.124323e-12, -2.356115e-11, -1.650269e-12, 
    -8.074985e-12, -7.087386e-13, 2.287143e-12, 5.874293e-12, 7.131629e-12, 
    1.014278e-11, -7.107724e-11, 1.484424e-12, 1.347344e-11, -1.573319e-11, 
    -2.118417e-12, -9.408385e-11, -8.508416e-12, -7.416481e-13, 4.751588e-12, 
    9.168999e-12, -8.777268e-12, -6.116774e-13, 6.242917e-12, 6.160739e-12, 
    -1.696043e-12, -9.126189e-12, -9.686563e-11, -5.219158e-13, 
    -2.347011e-14, -8.059886e-12, -9.98529e-12, -1.89862e-13, 6.29808e-12, 
    6.003864e-12, 7.698731e-12, 6.24889e-12, -6.879608e-12, -1.327627e-11, 
    5.006551e-12, -1.425227e-11, -1.680267e-11, -8.094525e-12, -6.55509e-12, 
    2.604006e-11, 4.043765e-13, 8.210099e-14, -2.122219e-12, -2.049819e-12, 
    8.898215e-12,
  -2.868428e-11, 8.169909e-12, 7.76168e-12, 5.019429e-12, 1.112532e-11, 
    1.234246e-11, 1.185482e-10, 1.168639e-10, -8.823475e-11, -5.185896e-11, 
    1.641687e-12, -1.015632e-11, -2.763345e-11, -2.346523e-11, -6.350254e-11, 
    5.06829e-12, -5.425327e-13, -9.75009e-12, -5.444797e-12, -3.006484e-12, 
    4.315437e-12, 4.343492e-11, 4.930178e-11, -3.798295e-12, 1.486478e-11, 
    -6.47693e-12, -4.676004e-11, 1.536227e-11, 5.365486e-12, 2.02266e-11, 
    3.186107e-11, -3.00221e-11, 3.567047e-11, -9.741319e-12, 3.887857e-11, 
    -3.3476e-11, -7.845824e-12, 2.335285e-12, 2.411593e-11, 3.097478e-12, 
    -2.382183e-12, 2.518763e-12, -1.497802e-12, -1.001097e-12, 1.036038e-11, 
    -6.070811e-12, -9.986456e-13, 5.54834e-14, -2.346945e-12, 5.61988e-13, 
    2.783468e-13, -1.242351e-11, -3.100742e-13, -1.101053e-12, 6.394885e-13, 
    1.801337e-13, -1.152123e-11, 6.151413e-12, -1.447165e-12, 5.059296e-11, 
    -1.616451e-11, 3.13749e-13, 3.376521e-12, -1.331624e-12, -5.831247e-12, 
    4.896805e-11, -3.139722e-11, 3.770084e-11, 3.809264e-11, -1.208145e-12, 
    -5.343026e-11, -1.749401e-11, -8.024248e-12, -1.294309e-11, 4.746315e-13, 
    -3.164247e-12, -6.619427e-13, 3.718692e-12, -4.785866e-13, 5.791922e-12, 
    4.373668e-12, -7.585952e-11, 8.307799e-13, 2.702316e-11, -1.911249e-11, 
    1.102196e-11, 1.965561e-11, -8.357204e-12, 1.032844e-12, 6.337375e-12, 
    2.084188e-11, -1.089018e-11, -7.672474e-13, 1.067023e-11, 3.549383e-12, 
    5.386624e-12, -8.839663e-12, 4.733158e-11, -5.014877e-13, -2.364464e-12, 
    -1.925882e-11, -2.210035e-11, 1.169939e-12, 6.81518e-12, -4.067191e-12, 
    -1.387956e-11, 7.882583e-13, 7.396417e-12, -2.166045e-12, 5.239031e-12, 
    -1.317557e-11, -1.68251e-11, -4.3755e-12, -2.520761e-12, 3.213563e-11, 
    2.754574e-13, 1.878775e-13, -8.596734e-13, 9.254923e-12, 6.966538e-12,
  -3.042167e-11, 3.980638e-11, 2.465583e-11, 4.015077e-11, 6.880962e-11, 
    1.346143e-10, 1.196778e-10, 6.71101e-11, -3.965761e-11, 1.083533e-11, 
    -1.385558e-12, -6.086176e-11, -9.158452e-12, 1.933498e-11, -5.481748e-11, 
    3.264322e-12, -2.876588e-13, -5.168532e-12, -5.742296e-12, 1.008726e-11, 
    1.189382e-11, 1.693579e-11, 4.830247e-11, -2.507328e-12, 6.779155e-11, 
    -7.189316e-11, -1.432388e-11, 3.048006e-11, 6.775913e-12, 2.601741e-11, 
    -3.642375e-11, 2.058287e-11, -6.315437e-11, -3.244072e-13, 1.107225e-11, 
    5.871437e-11, -2.245226e-12, 1.062817e-12, 4.936052e-13, 2.889289e-12, 
    -1.367253e-11, 1.247891e-12, -3.733347e-12, -3.836546e-12, -5.33884e-12, 
    -2.784661e-11, -2.364331e-12, 1.206035e-12, -7.812373e-12, -5.125067e-13, 
    3.524042e-12, -2.754996e-11, -2.247935e-12, -3.639311e-13, 1.319739e-12, 
    4.194423e-13, 3.962741e-11, 4.065192e-13, -1.598255e-12, 9.582302e-11, 
    1.310152e-11, -3.539613e-12, -2.230771e-11, -2.826583e-12, -4.882717e-12, 
    9.210743e-11, -1.863401e-10, 2.097456e-11, 1.144818e-11, 2.575717e-13, 
    -9.205969e-12, -2.41942e-11, -1.552758e-11, -4.116019e-11, -2.084999e-12, 
    4.602985e-13, -3.839706e-13, 6.330214e-12, -1.332701e-12, 6.456835e-12, 
    4.247713e-13, -4.224201e-11, -3.657075e-13, 6.445733e-12, 4.440892e-16, 
    4.147815e-11, -3.433454e-11, -1.382294e-11, 1.016829e-12, 6.403322e-12, 
    2.497691e-11, -1.551466e-11, -1.305678e-12, 8.606649e-12, -5.423972e-11, 
    3.297296e-12, -2.47713e-12, -7.618128e-12, -8.987255e-12, -3.007372e-12, 
    -1.97522e-11, -1.367796e-11, 2.901165e-12, 6.164513e-14, 1.90612e-11, 
    -2.971556e-11, 1.377343e-11, 2.49516e-11, 1.428213e-11, 8.572698e-12, 
    -8.447465e-12, -7.470691e-12, 2.977174e-12, 5.192735e-12, 3.378031e-11, 
    1.833422e-13, 1.889044e-13, 1.213488e-12, 1.435131e-11, 8.926415e-12,
  9.402656e-11, -9.684031e-12, 4.659495e-11, 9.210477e-11, 1.692839e-10, 
    1.70115e-10, 8.676504e-11, -8.761325e-11, -1.663403e-10, 2.273004e-10, 
    1.305547e-10, -1.052392e-10, 2.880962e-11, 3.297629e-11, 3.399947e-12, 
    9.25926e-13, -4.579448e-13, -4.96847e-12, -4.926615e-12, -2.866152e-12, 
    2.664069e-11, 2.324496e-11, 3.613843e-11, -1.226801e-10, 9.132251e-11, 
    -5.716205e-11, 8.940115e-11, 6.528511e-11, 3.766965e-11, 5.173906e-11, 
    -2.900902e-11, 1.570295e-10, -2.554794e-10, 3.503065e-11, 3.662182e-12, 
    6.708611e-11, -1.871459e-12, 3.005929e-13, -3.807421e-11, 2.326428e-12, 
    -1.253193e-11, -7.530865e-12, -6.528778e-12, -4.90729e-12, -1.427769e-11, 
    -7.696288e-11, -3.953948e-12, -4.50362e-13, -1.576703e-11, -1.640785e-12, 
    3.615858e-12, -8.816503e-12, -4.491074e-13, 5.402345e-13, 7.200518e-13, 
    6.140644e-13, 1.259726e-11, -2.636647e-12, -1.370735e-11, 2.924519e-11, 
    3.902345e-11, -1.899481e-11, -5.089573e-11, -6.534728e-12, -3.508838e-12, 
    8.440781e-11, 4.734804e-10, 1.932654e-11, 4.656941e-11, -2.69289e-11, 
    1.980816e-11, -5.314083e-11, 8.982015e-11, -1.076279e-10, -2.194034e-11, 
    2.946532e-13, -1.98036e-13, 5.598189e-12, -1.875533e-12, 2.809308e-12, 
    -1.208367e-12, -7.208018e-12, -2.655209e-12, -2.077849e-11, 2.338463e-11, 
    9.046852e-11, 6.605716e-11, -1.720579e-11, 8.645896e-13, 4.426237e-12, 
    1.429412e-11, -2.686202e-11, -1.885991e-12, 1.565259e-12, -7.767342e-11, 
    8.610757e-12, 4.488321e-12, 7.34568e-12, -1.779998e-11, -2.585798e-12, 
    -1.518585e-11, -1.054762e-11, 3.631234e-12, -3.946427e-13, 3.656364e-11, 
    -3.138112e-11, 1.632694e-11, 3.622258e-11, 1.635936e-11, 9.247492e-12, 
    -1.272094e-11, 3.599343e-12, 4.301892e-12, -1.159517e-12, 3.319567e-11, 
    1.939338e-13, -2.969569e-13, 9.848095e-13, 8.984383e-12, 6.523893e-12,
  1.518694e-10, -3.69933e-11, 6.078227e-11, 1.429978e-10, 1.785281e-10, 
    1.63572e-10, -1.118727e-11, -1.709031e-10, -9.810308e-11, 5.933323e-10, 
    -2.342035e-10, -2.941669e-11, 1.765892e-10, 3.047584e-11, -4.807021e-11, 
    -6.596057e-13, -1.38245e-13, -1.007372e-11, -4.830025e-12, -1.314748e-11, 
    6.257883e-12, 1.556155e-11, 7.298273e-11, -2.585521e-10, 5.980527e-11, 
    -3.145639e-11, 3.485678e-11, 1.415812e-10, 2.244183e-11, 1.110323e-10, 
    5.729883e-11, 1.107801e-10, 1.336786e-10, 6.686629e-11, -2.409473e-11, 
    -6.226797e-12, 2.159295e-12, 1.24234e-13, 2.787703e-11, -8.278711e-13, 
    7.882538e-12, -1.912359e-11, -7.996381e-12, 1.21525e-12, 2.570988e-11, 
    -3.547052e-11, -4.692469e-12, -3.510192e-12, -3.07161e-11, -2.111783e-12, 
    1.106476e-11, -1.775091e-11, 1.356515e-12, -3.126255e-12, 5.104805e-14, 
    -4.818368e-14, 1.131821e-10, -4.392664e-12, -2.210068e-11, 2.305905e-11, 
    4.144307e-11, -2.245648e-11, -5.227974e-11, -1.140106e-11, -6.963186e-12, 
    9.647327e-11, 1.874834e-11, 1.564044e-10, -9.104495e-12, -9.533196e-11, 
    9.751244e-11, -9.840595e-11, 1.7613e-10, -9.357648e-11, -4.445302e-11, 
    6.639134e-14, 8.715251e-15, 1.576628e-12, -6.610046e-13, -1.107492e-11, 
    -3.602452e-12, 2.875276e-11, -4.548362e-12, 1.486702e-10, -1.772398e-10, 
    1.585156e-10, 2.018614e-10, -1.776113e-11, 6.006723e-13, 1.275202e-12, 
    -6.826317e-12, -2.03928e-11, -1.720069e-12, -1.948064e-11, -7.774381e-11, 
    9.376455e-12, 9.390044e-12, 1.815548e-11, -1.251199e-11, -2.412426e-12, 
    -3.059175e-11, -7.280399e-12, 2.903261e-12, 8.19067e-14, 5.760836e-11, 
    -1.983547e-11, 5.52165e-11, 4.884559e-11, 4.664935e-12, 7.730039e-12, 
    -1.168687e-11, 1.023071e-11, 1.111444e-11, -1.211053e-11, 4.356138e-11, 
    2.627676e-13, -1.875222e-12, -6.566969e-14, 5.192902e-12, 1.238321e-11,
  1.162523e-10, -1.517941e-11, 6.366774e-11, 1.288645e-10, 1.704312e-10, 
    1.224323e-10, -1.388485e-10, -9.84044e-11, 1.891154e-11, 4.79806e-10, 
    -7.28515e-11, -2.750289e-11, 8.700285e-11, -1.786082e-11, -1.649441e-10, 
    -2.83098e-12, -8.138379e-13, -1.568612e-11, -8.637868e-12, -8.523404e-12, 
    2.571721e-12, -4.654499e-12, 2.494294e-10, 1.664477e-10, 1.035483e-11, 
    -1.503353e-10, 3.160983e-11, 2.109277e-10, 3.275735e-11, 1.613567e-10, 
    1.2473e-10, 1.068412e-10, 1.392881e-10, 1.237068e-10, -1.674794e-11, 
    -7.524203e-12, 3.579181e-12, 1.103562e-13, -3.05449e-11, -8.014389e-12, 
    7.301937e-11, -3.631451e-11, -2.045253e-12, 5.878964e-12, 9.003776e-11, 
    -1.289711e-10, -9.945822e-12, -4.279022e-12, -5.140697e-11, 
    -6.709633e-13, 1.58954e-11, -4.391465e-11, -6.027268e-12, -1.129168e-11, 
    5.705436e-13, -4.214407e-13, -8.476375e-11, -1.052376e-11, -2.412692e-11, 
    8.852374e-11, 3.268097e-11, -1.073852e-11, -1.746603e-12, -1.201625e-11, 
    -8.111112e-12, 1.319793e-10, 4.460676e-10, 2.24889e-10, 5.928991e-11, 
    -2.041705e-10, 1.562701e-10, -1.02681e-10, 5.815837e-11, 3.999512e-11, 
    -6.20056e-11, -2.436717e-12, 2.200462e-13, 5.441203e-12, 2.606049e-12, 
    -2.465894e-11, -8.716139e-12, 6.141476e-11, -9.132251e-12, 3.731357e-10, 
    -1.235114e-10, 1.536136e-10, 4.902039e-10, -3.203171e-11, -1.855738e-13, 
    -1.065814e-12, -3.478773e-11, -1.646372e-11, -1.026956e-12, 
    -3.008935e-11, -3.536682e-11, -1.115481e-11, 1.669411e-11, -6.948664e-12, 
    -4.971579e-12, -1.429168e-12, -4.356915e-11, 1.411626e-11, 6.10012e-13, 
    1.352918e-12, 2.060174e-11, -2.82574e-12, 1.019376e-10, 2.605871e-11, 
    -2.913669e-12, 7.6672e-12, 9.738876e-13, 2.545564e-11, 1.814238e-11, 
    7.621015e-12, 6.091083e-11, 9.281464e-14, -3.529399e-12, -4.493073e-13, 
    3.872791e-12, 4.35576e-11,
  6.592771e-11, 2.714096e-11, 4.123635e-11, 9.935874e-11, 1.774865e-10, 
    3.427658e-11, -2.002114e-10, 1.029434e-10, 1.610854e-10, 7.748469e-12, 
    8.490986e-13, -9.815082e-11, -3.037748e-11, -7.40723e-11, -2.478018e-10, 
    -6.413003e-12, -1.961098e-12, -1.450129e-11, -1.088729e-11, 5.369927e-12, 
    2.944844e-11, -2.266987e-11, 2.437783e-10, 9.139267e-10, -1.724558e-10, 
    -2.610392e-10, 1.101093e-10, 3.075158e-10, 8.145129e-11, 1.809521e-10, 
    -4.949641e-11, 3.058105e-10, -9.628565e-11, 2.129266e-10, -6.027179e-12, 
    2.309921e-10, 5.615064e-13, -4.996004e-14, -2.514664e-10, -1.772449e-11, 
    1.997815e-10, -1.149676e-10, 1.111866e-11, 6.59961e-12, 6.392042e-11, 
    -3.758558e-10, -2.909051e-11, -7.491785e-12, -6.50946e-11, 6.004974e-12, 
    2.062817e-11, -3.303668e-11, -2.334009e-11, -1.397247e-11, 1.274136e-12, 
    -5.062617e-13, -2.267537e-10, -2.770619e-11, -3.790639e-11, 2.633191e-10, 
    4.355982e-11, -3.5147e-11, 4.934186e-11, -8.460077e-12, -1.909939e-12, 
    1.793925e-10, 1.00643e-09, -1.748202e-10, 2.244569e-10, -3.343068e-10, 
    1.544009e-10, -2.364455e-10, -2.80215e-10, 1.10477e-10, -6.049401e-11, 
    -1.109868e-11, 2.196021e-13, 2.25886e-11, 8.980194e-12, -2.979306e-11, 
    -1.583356e-11, 8.248575e-11, -1.15179e-11, 5.807834e-10, -3.307576e-12, 
    8.075673e-11, 7.046701e-10, -4.816059e-11, -3.973488e-13, -1.483258e-12, 
    -9.901058e-11, -1.918963e-11, -3.863576e-13, -2.843486e-11, 8.686385e-13, 
    -5.856134e-11, 2.958984e-11, 2.23519e-11, -1.294076e-11, -2.163603e-13, 
    -7.272938e-11, 4.62147e-11, -1.199152e-12, 3.41116e-12, -6.068035e-12, 
    -9.424816e-11, 4.613376e-11, -5.825562e-11, 5.265122e-12, 3.568701e-12, 
    1.884715e-12, 5.424816e-11, 3.722178e-11, 4.208722e-11, 8.51994e-11, 
    6.412648e-14, -3.319789e-12, -2.691181e-13, 2.98539e-12, 5.793765e-11,
  5.788436e-11, 1.06775e-10, 3.646861e-12, 6.849632e-11, 1.704397e-10, 
    1.14575e-12, -1.922587e-10, 3.530864e-10, 4.21938e-10, -2.670379e-10, 
    -2.195399e-11, -1.141949e-10, -7.968026e-11, -1.358718e-10, 
    -3.042651e-10, -1.260894e-11, -3.235101e-12, -3.453238e-12, 
    -1.074629e-11, 2.450662e-11, 5.47935e-11, -3.645262e-11, 7.743495e-11, 
    1.29611e-09, -5.695142e-10, -3.15822e-10, 2.250538e-10, 3.527418e-10, 
    3.307594e-10, 1.081126e-10, 3.579821e-10, 3.558398e-10, -3.661906e-10, 
    1.747331e-10, 5.529088e-11, -7.003997e-11, -2.149925e-12, -3.506084e-13, 
    -2.094378e-10, -3.044729e-11, 2.563983e-10, -2.390728e-10, 2.11231e-11, 
    5.420192e-12, -1.24933e-10, -5.013092e-10, -7.266721e-11, -2.154765e-11, 
    -7.31557e-11, 1.195666e-11, 2.344813e-11, 2.999734e-11, -2.824212e-11, 
    -8.408563e-12, 1.323164e-12, -1.047162e-12, -6.09468e-10, -6.891145e-11, 
    -8.294876e-11, 3.921492e-10, 8.65974e-11, -1.327098e-10, 9.500489e-11, 
    -6.22471e-12, 3.012346e-12, 2.018687e-10, 3.352095e-09, 2.115623e-10, 
    3.414975e-10, -4.389324e-10, 2.107896e-10, -1.880185e-10, 5.842082e-11, 
    6.464163e-11, -4.70882e-11, -2.267342e-11, 1.310063e-14, 4.928502e-11, 
    1.885634e-11, -1.314504e-12, -3.148237e-11, 9.90442e-11, -1.389733e-11, 
    2.036558e-10, -8.602541e-11, 1.046949e-10, 1.275714e-09, -5.799983e-11, 
    2.027795e-12, -8.348877e-14, -3.00405e-10, 9.525358e-11, 4.982681e-13, 
    -4.967813e-11, -9.195489e-11, -1.217618e-10, 5.79135e-11, 1.375948e-10, 
    -3.874057e-11, -3.28626e-13, -1.00826e-11, 8.53968e-11, -3.608447e-12, 
    4.046319e-12, 2.776623e-11, -3.345431e-10, -1.280434e-10, -1.595826e-10, 
    -2.120792e-11, 8.331114e-12, 4.005685e-12, 8.10676e-11, 7.790391e-11, 
    7.476686e-11, 1.067306e-10, 1.124434e-13, -1.777023e-12, 8.382184e-13, 
    4.698464e-13, 3.59357e-11,
  7.366197e-11, 1.707772e-10, 9.503509e-13, 5.298695e-11, 2.400178e-10, 
    1.383214e-10, -1.676081e-10, 5.448477e-10, 1.368626e-09, 1.338858e-10, 
    -1.017852e-10, 2.197762e-10, 3.446115e-10, -1.576534e-10, -3.585026e-10, 
    -1.873026e-11, -3.92788e-12, 1.578293e-11, -7.503997e-12, 4.387601e-11, 
    6.181722e-11, -4.982859e-11, 6.067147e-11, 1.249466e-09, -5.400462e-10, 
    -2.791687e-10, 3.572396e-10, 1.137712e-09, 8.905463e-10, 1.831033e-10, 
    8.070629e-10, 4.177707e-10, -4.494449e-10, -3.919176e-11, -5.736744e-11, 
    6.77769e-11, 6.267697e-12, 3.708145e-14, 9.535484e-11, -5.225189e-11, 
    2.590067e-10, -2.886598e-10, 2.090195e-11, -2.275791e-12, -2.604796e-10, 
    -9.977708e-10, -1.475513e-10, -5.086065e-11, -7.617373e-11, 
    -5.310974e-12, 1.383449e-11, 2.487592e-10, -1.928484e-11, -1.987033e-12, 
    4.56124e-13, -2.481571e-12, -1.068454e-09, -1.585027e-10, -2.733447e-10, 
    2.920069e-10, 1.780567e-10, -2.651959e-10, 1.113616e-10, 1.979217e-12, 
    4.324719e-12, 5.803891e-11, 2.491433e-09, 5.244445e-10, 5.098926e-10, 
    -5.07848e-10, 6.6807e-10, 6.110845e-11, -1.415453e-09, -4.443024e-11, 
    -5.02137e-11, -3.376144e-11, 2.68674e-13, 7.791146e-11, 2.919163e-11, 
    -1.016947e-10, -5.87832e-11, 1.116311e-10, -1.826628e-11, 7.398793e-10, 
    4.336531e-10, -1.788365e-10, 2.04877e-09, -5.403855e-11, 1.08642e-11, 
    8.646417e-12, -4.049792e-10, 2.172026e-10, 1.502798e-12, -7.132925e-11, 
    -1.139533e-11, -1.678082e-10, 9.962449e-11, 2.454801e-10, -7.416112e-11, 
    3.176481e-12, 1.267679e-10, 1.75398e-10, -1.103528e-11, 1.131983e-12, 
    1.790532e-10, -5.55783e-10, -1.554241e-10, -2.391864e-10, -3.017444e-10, 
    -5.077361e-11, -9.618972e-12, 1.134524e-10, 1.371898e-10, 9.937828e-11, 
    1.018172e-10, 1.601208e-12, -4.563017e-13, 3.204714e-12, -4.539258e-12, 
    -2.748024e-11,
  8.126122e-11, 7.510081e-11, -7.492673e-11, 4.525447e-11, 4.050875e-10, 
    4.411582e-10, -3.516121e-11, 3.852385e-10, 2.320267e-09, 1.503651e-09, 
    -2.31914e-10, 6.50882e-10, 8.613874e-10, -1.386766e-10, -3.781579e-10, 
    -1.190692e-11, -3.554845e-12, 3.873879e-11, -2.434053e-12, 5.917045e-11, 
    5.929124e-11, -5.653789e-11, 2.272564e-10, 7.683099e-10, -9.346834e-11, 
    9.993428e-11, 3.451603e-10, 1.391403e-09, 1.364047e-09, 3.306759e-10, 
    1.607301e-09, 5.21041e-11, -1.695355e-11, -4.606093e-11, -9.321965e-11, 
    4.862919e-10, 2.237108e-11, 4.119372e-12, 5.521912e-10, -9.96419e-11, 
    -5.161382e-12, -2.542926e-10, -5.666578e-13, -2.178213e-11, 
    -4.955325e-10, -3.969411e-10, -2.487415e-10, -9.894574e-11, 
    -9.081518e-11, -4.711898e-11, 6.199086e-11, 5.075655e-10, -4.746284e-11, 
    3.540066e-11, 9.95648e-14, -4.069634e-12, -2.153662e-09, -3.214925e-10, 
    -3.804978e-10, 2.678751e-10, 3.071108e-10, -3.577441e-10, 1.407763e-10, 
    1.761364e-11, 1.033698e-11, -2.802736e-10, 1.473772e-10, 2.232714e-09, 
    4.190071e-10, -6.764829e-10, 1.352131e-09, 5.592327e-11, 1.159187e-09, 
    -1.046629e-10, -9.204512e-11, -4.096279e-11, 1.07736e-12, 6.484147e-11, 
    2.440759e-11, -6.668017e-10, -8.324186e-11, 1.333341e-10, -2.368772e-11, 
    8.368559e-10, 5.374794e-10, -6.436061e-10, 2.04216e-09, -4.51692e-11, 
    3.657524e-11, 2.878231e-11, -7.43988e-10, -1.040739e-10, 2.202682e-12, 
    -2.198384e-11, 2.34408e-10, -3.261111e-10, 1.687809e-10, 2.518163e-10, 
    -1.037606e-10, -5.683631e-12, 7.823431e-11, 3.408385e-10, -2.834888e-11, 
    -3.120393e-12, 4.333707e-10, -5.120278e-10, -1.942944e-10, 1.754898e-10, 
    -5.881589e-10, -2.275549e-10, -3.604228e-11, 1.309672e-10, 1.892104e-10, 
    1.471818e-10, 5.605472e-11, 4.17586e-12, 8.864021e-13, 5.746847e-12, 
    -6.969536e-12, -1.121805e-10,
  4.974154e-11, 1.134559e-10, -7.462475e-11, -2.061462e-10, 2.0027e-10, 
    5.56593e-10, 4.562715e-10, -4.676437e-11, 9.023218e-10, 1.995399e-09, 
    -7.084644e-10, 7.968985e-10, -1.631665e-09, -9.441337e-11, -2.914895e-10, 
    4.276828e-11, -2.938165e-11, 6.461676e-11, 1.442135e-11, 6.549428e-11, 
    4.961365e-11, -2.471623e-11, 2.271072e-10, 2.486509e-10, -8.766143e-10, 
    3.580958e-10, 8.643646e-10, 1.702102e-09, 1.182496e-09, 3.448015e-10, 
    3.948667e-09, 5.024781e-10, -2.435137e-10, 2.288765e-10, -1.075939e-10, 
    1.012477e-09, 1.931966e-11, 1.029576e-11, 7.181349e-10, -1.923816e-10, 
    2.140162e-10, -2.2089e-10, -3.370282e-11, -8.26833e-11, -1.143821e-09, 
    -5.403358e-10, -3.92923e-10, -1.82121e-10, -1.996447e-10, 4.363176e-12, 
    3.755387e-10, 1.748894e-10, -6.972343e-11, 8.444303e-11, 7.366374e-12, 
    -3.641532e-12, -3.387203e-09, -5.640928e-10, -4.34319e-11, 4.252572e-10, 
    4.616787e-10, -4.210641e-10, 7.311129e-11, 2.434248e-11, 3.57538e-11, 
    -5.550937e-10, 7.084289e-10, -3.748362e-10, 2.738947e-09, -7.477432e-10, 
    9.98984e-10, -1.89825e-10, 1.28551e-09, -8.299175e-10, -1.965418e-10, 
    -3.634781e-11, 1.159073e-12, -1.293188e-11, 4.156675e-14, -5.92717e-10, 
    -9.909584e-11, 1.607926e-10, -2.881606e-11, 1.884583e-09, 4.565397e-09, 
    5.046878e-10, 1.248015e-09, -4.140688e-11, 8.750223e-11, 4.554934e-11, 
    -1.849909e-09, -4.242786e-10, -3.009148e-12, 2.913652e-11, 1.317677e-09, 
    -8.847345e-10, 2.565066e-10, 4.613092e-10, -1.311342e-10, -2.890559e-11, 
    -1.169873e-10, 5.428342e-10, -5.190159e-11, 2.938982e-12, 6.717791e-10, 
    -1.932854e-10, -3.745591e-10, 3.391882e-10, -1.100187e-09, -2.76696e-10, 
    -1.064144e-10, 3.806022e-11, 2.328839e-10, 2.263896e-10, -4.654055e-13, 
    6.131273e-12, 4.908074e-12, 6.808776e-12, -1.100675e-11, -1.974918e-10,
  7.81526e-11, 8.279954e-11, 3.511644e-10, 4.905942e-10, -6.910739e-11, 
    -4.926193e-11, 7.049579e-10, 6.904344e-11, -7.801759e-11, 1.050722e-09, 
    -7.369039e-11, 6.792504e-10, -8.757866e-10, -2.33058e-11, -1.875335e-10, 
    -2.225285e-10, -1.437975e-10, 7.699796e-11, 3.729195e-11, 3.985434e-11, 
    4.122569e-11, 5.28857e-11, 1.983551e-10, 2.203606e-10, -5.732872e-10, 
    -1.996199e-09, 4.100613e-10, 4.204388e-09, 9.045422e-10, -9.541878e-11, 
    8.014489e-09, 1.539831e-09, 5.501093e-10, 1.021121e-10, -2.346141e-10, 
    1.074945e-09, -5.261001e-11, 1.501821e-11, -5.850467e-10, -3.028781e-10, 
    5.864038e-10, -2.890133e-10, -4.496492e-11, -1.945115e-10, -1.992802e-09, 
    -6.026113e-10, -5.831566e-10, -2.858727e-10, -4.866251e-10, 1.43149e-10, 
    9.761481e-10, -6.642722e-10, -1.107061e-10, 1.143363e-10, 2.797904e-11, 
    1.488587e-12, -3.839972e-09, -8.783737e-10, -5.435176e-10, 8.424736e-10, 
    5.53726e-10, -4.746781e-10, -1.16458e-11, 1.689955e-11, 4.521468e-11, 
    -5.139427e-10, 4.613518e-09, 8.851941e-10, 7.890577e-10, -1.138545e-09, 
    -6.330723e-10, -8.957315e-10, 9.274004e-10, -1.263629e-09, -3.162846e-10, 
    -9.15179e-12, 1.90159e-12, -1.685976e-10, -1.816591e-11, 1.271729e-10, 
    -9.815082e-11, 1.917194e-10, -3.61382e-11, 3.405837e-09, 2.176392e-09, 
    2.004249e-09, 1.173461e-10, -3.211653e-11, 1.304803e-10, 4.227019e-11, 
    2.958416e-10, -3.308614e-10, -1.545253e-11, -1.294745e-09, 3.85036e-09, 
    -1.710204e-09, 3.621281e-10, 1.017369e-09, -1.58515e-10, -6.205454e-11, 
    -8.279244e-11, 6.984178e-10, -9.268364e-11, 2.692069e-11, 5.499246e-10, 
    -3.235101e-11, -2.276366e-10, -3.489191e-10, -3.761116e-10, 3.768292e-10, 
    -1.656204e-10, -1.913705e-10, 1.581455e-10, 3.346301e-10, -8.91589e-11, 
    9.705303e-12, 1.090683e-11, 8.033352e-12, -1.267386e-11, -2.938378e-10,
  1.582769e-10, 2.634657e-10, 2.392266e-09, 4.801333e-09, -4.240412e-10, 
    -2.120547e-09, -6.142642e-12, 6.026646e-10, -3.490932e-10, -1.624052e-10, 
    1.911467e-10, 5.686012e-10, -1.549445e-10, 8.465051e-11, -5.517364e-12, 
    -4.60016e-10, -3.372308e-11, -4.139267e-11, 6.191314e-11, -3.744915e-11, 
    4.852652e-11, 1.434977e-10, 2.044906e-10, 9.433556e-10, 2.717837e-09, 
    -4.768285e-09, -8.566765e-10, 7.549087e-09, 1.495618e-09, -5.80048e-10, 
    5.43471e-09, 6.88058e-09, 6.904852e-09, -1.041773e-09, -5.982663e-10, 
    2.976144e-10, -1.619945e-10, 2.345857e-11, 3.4977e-09, -3.558391e-10, 
    7.947612e-10, -5.546674e-10, -4.131451e-11, -2.393967e-10, -2.840597e-09, 
    -3.078391e-10, -7.851177e-10, -3.146461e-10, -5.659878e-10, 1.180469e-10, 
    1.626971e-09, -5.053558e-10, -1.883628e-10, 1.093376e-10, 3.111751e-11, 
    1.122302e-11, -2.844846e-09, -1.238853e-09, -1.632544e-09, -8.645706e-10, 
    4.973479e-10, -5.678551e-10, -4.161116e-10, -3.994742e-11, 9.671198e-12, 
    -7.313652e-10, 1.563645e-09, -1.076902e-09, 2.038902e-11, -2.163265e-09, 
    -1.955957e-09, -1.043762e-09, 7.462937e-10, -7.057714e-10, -3.583416e-10, 
    1.628209e-11, 4.517275e-12, -4.163176e-10, -1.711129e-11, 2.035669e-10, 
    -8.074252e-11, 1.886949e-10, -5.776357e-11, 4.668063e-09, 2.980581e-09, 
    8.475887e-10, -1.35012e-09, -2.778577e-11, 1.630627e-10, 1.891003e-10, 
    3.452453e-09, 1.113129e-10, -2.196288e-11, -6.250353e-09, 2.493277e-09, 
    -2.44049e-09, 4.698727e-10, 1.422674e-09, -1.645226e-10, -7.105498e-11, 
    3.855938e-10, 7.081677e-10, -1.966995e-10, 5.726353e-11, 2.196963e-10, 
    4.251568e-10, -1.783782e-10, -3.027555e-09, -2.777742e-09, 2.415273e-09, 
    -1.203126e-10, -3.292406e-10, -2.791367e-11, 8.344294e-10, -2.776552e-10, 
    1.440199e-11, 1.853806e-11, 1.72431e-11, -1.313616e-11, -4.134542e-10,
  1.16561e-10, 3.132886e-09, 8.445813e-09, 3.649365e-09, -5.832472e-09, 
    -5.384347e-09, -3.885472e-09, 5.945715e-10, 4.786571e-11, 2.848175e-10, 
    1.10936e-09, 7.630128e-10, 2.264205e-09, 1.46489e-10, 1.103366e-10, 
    1.451761e-10, -8.925048e-10, -6.162857e-10, 3.857359e-11, -7.736034e-11, 
    7.667111e-11, 2.462919e-10, 2.016698e-10, 1.213127e-09, 3.60281e-09, 
    -4.712426e-10, -6.164314e-11, 9.087618e-09, -2.872962e-09, -1.572584e-09, 
    2.485866e-09, 1.088961e-08, 6.415679e-09, -2.698709e-09, -1.343334e-09, 
    -8.603784e-10, -1.644985e-10, 2.277289e-11, 9.027662e-09, -2.643482e-10, 
    6.077478e-10, -1.166409e-09, 1.124185e-10, -2.951617e-11, -4.351559e-09, 
    6.709406e-10, -1.609809e-09, 1.035261e-11, 2.419519e-10, 6.874057e-11, 
    1.378291e-09, -2.426752e-10, -1.163578e-10, 8.283862e-11, 1.488623e-11, 
    1.693579e-11, -4.393012e-09, -2.200917e-09, -2.841731e-09, 4.977863e-09, 
    3.777849e-10, -7.368861e-10, -1.184755e-09, -9.347012e-10, 1.123351e-12, 
    -1.605425e-09, 5.271978e-10, -2.604533e-09, -1.129759e-09, -2.619132e-09, 
    -1.728079e-09, -1.683485e-09, -5.533387e-10, -2.082015e-09, 
    -2.769731e-10, 1.650236e-11, 1.159073e-11, -8.720527e-10, -1.196849e-10, 
    4.415917e-10, 5.830003e-12, 1.913499e-10, -1.070326e-10, 6.231122e-09, 
    -2.859046e-10, -1.047304e-10, -3.434121e-09, -2.210854e-11, 2.28088e-10, 
    5.478533e-10, 7.338119e-09, -2.473534e-10, -2.182787e-11, -6.073268e-09, 
    7.335252e-10, -3.999147e-09, 5.482896e-10, 2.291959e-09, -1.308642e-10, 
    -8.386607e-11, 1.245073e-09, 4.828458e-10, -3.979848e-10, 9.941736e-11, 
    1.089266e-09, 1.058034e-10, -9.735821e-10, -2.877339e-09, 6.893437e-10, 
    4.703839e-09, -1.261746e-10, -2.244995e-10, -1.692335e-10, 9.757493e-10, 
    -4.372644e-10, 1.848335e-11, 2.150102e-11, 4.177014e-11, -2.361578e-11, 
    -5.57332e-10,
  6.945555e-12, 7.656421e-09, 1.163574e-08, 1.228404e-08, 2.59659e-09, 
    -6.542809e-09, -9.394501e-09, -8.814034e-10, 1.119854e-09, 1.113914e-09, 
    2.854488e-09, 1.756842e-09, 6.550742e-10, -1.36982e-10, -1.964118e-10, 
    2.347811e-11, -1.617446e-09, -4.646985e-10, 1.783462e-11, -8.062173e-11, 
    1.290168e-10, 4.207941e-10, 6.080469e-11, 7.141061e-10, 1.008811e-09, 
    1.525688e-09, 3.037012e-09, 5.966069e-09, 4.752462e-09, -3.355996e-09, 
    1.200998e-09, 1.1158e-08, 4.238625e-09, -1.268564e-09, -2.197783e-09, 
    -3.622848e-09, -7.790746e-11, 1.659473e-11, -1.021379e-08, -2.468177e-10, 
    5.367773e-10, -1.902908e-09, 1.975486e-10, -1.569891e-10, -6.772058e-09, 
    1.187839e-09, -5.211692e-09, 1.431779e-10, 8.956015e-10, 7.401901e-11, 
    5.578293e-10, -2.971667e-10, 2.765645e-11, 6.857519e-11, -4.178702e-12, 
    4.543921e-12, -4.726434e-09, -5.68353e-09, -8.300805e-09, 1.968846e-09, 
    4.614655e-10, -1.116536e-09, -1.621419e-09, -3.156499e-09, 1.450541e-09, 
    -1.631168e-09, 1.088487e-08, -4.058382e-09, -1.243382e-09, -2.384141e-09, 
    -1.943324e-09, -1.434621e-10, -4.042068e-09, -4.851547e-09, 8.402808e-11, 
    7.798207e-12, 2.410516e-11, -1.67832e-09, -2.940453e-10, 4.149609e-09, 
    1.700577e-10, 2.625377e-10, -1.640963e-10, 7.722047e-09, -2.501896e-09, 
    7.381793e-10, -5.215487e-09, 1.680789e-11, 1.658655e-10, 6.421423e-10, 
    1.092245e-08, -9.284641e-10, -2.328093e-11, 2.241613e-09, 2.696492e-09, 
    -7.085877e-09, 6.204679e-10, 4.261619e-09, -1.031317e-10, -7.318661e-11, 
    -1.348884e-09, 1.591793e-11, -6.514789e-10, 1.194955e-10, 1.193524e-09, 
    -2.114753e-10, -7.860379e-11, 7.009469e-10, 1.121617e-09, 4.242917e-09, 
    2.222684e-10, -2.1247e-10, -3.089333e-10, 7.146177e-10, -5.379555e-10, 
    4.328839e-11, 8.668621e-12, 7.204903e-11, -5.898038e-11, -7.712693e-10,
  1.399769e-10, 8.524552e-09, 9.153695e-09, 8.897558e-09, 6.102056e-09, 
    4.69052e-09, -7.548891e-09, -6.322409e-09, 8.076029e-10, 1.226169e-09, 
    4.606619e-09, -2.758043e-10, 2.614513e-10, 1.203063e-09, -1.125528e-09, 
    5.88082e-10, -2.893967e-09, 8.132304e-10, -5.267609e-11, 2.818297e-10, 
    1.518288e-10, 7.491394e-10, -8.677148e-11, 2.119407e-10, -3.910259e-10, 
    2.509438e-09, 6.488563e-09, 7.090108e-09, 1.651671e-08, -6.590454e-09, 
    4.135984e-09, 1.313742e-08, 1.042537e-09, 9.529515e-10, -1.431374e-09, 
    -6.502518e-09, -2.090417e-11, 3.144152e-12, -2.810222e-08, -4.428471e-10, 
    6.867481e-10, -2.023768e-09, -2.360707e-10, -5.225975e-10, -7.58746e-09, 
    2.904102e-09, -1.434478e-08, -1.906599e-10, 1.038154e-09, 8.626699e-11, 
    -7.231904e-11, -9.910082e-10, 3.200455e-10, 7.753442e-11, -1.177298e-11, 
    -3.82272e-11, -4.463885e-09, -1.166439e-08, -1.591538e-08, 5.966108e-10, 
    6.497487e-10, -1.695753e-09, -1.633595e-09, -5.820499e-09, 3.047063e-09, 
    -1.062091e-09, 1.072539e-08, -5.581938e-09, -9.552309e-09, -6.969003e-11, 
    -1.009965e-09, 9.539463e-10, -2.984507e-09, -3.258435e-09, 9.566974e-10, 
    4.158096e-11, 2.651035e-11, -2.170545e-09, -3.070156e-10, 6.675918e-09, 
    3.07125e-10, 4.60625e-10, -1.779625e-10, 9.562854e-09, -7.273229e-09, 
    2.297384e-09, -5.54482e-09, 1.235492e-10, -8.822942e-11, 1.051603e-12, 
    1.104215e-08, -1.0186e-09, -8.171241e-12, 3.84339e-09, 2.890289e-09, 
    -1.013334e-08, 5.736638e-10, 5.38779e-09, -8.157031e-11, -4.478125e-11, 
    -3.113996e-09, -1.151683e-10, -9.93797e-10, 1.043592e-10, 7.593997e-10, 
    5.096297e-10, 1.921222e-09, 2.578929e-09, -3.707925e-09, 4.915194e-09, 
    1.069509e-10, -2.374918e-10, -5.906315e-10, -1.707861e-10, -7.242136e-10, 
    8.203358e-11, 8.366641e-12, 8.71605e-11, -1.128697e-10, -9.688108e-10,
  2.114291e-10, 5.389012e-09, 6.13727e-09, 2.52183e-09, 4.816229e-09, 
    3.444683e-09, -3.117862e-11, -1.310426e-08, -1.561887e-09, 1.567713e-09, 
    3.298709e-09, -4.485884e-09, 4.01883e-10, -3.582841e-10, -1.582464e-09, 
    -4.93642e-10, -5.814897e-09, 1.439957e-09, -5.939427e-11, 6.600942e-10, 
    -2.854108e-10, 1.102705e-09, 9.271162e-11, 1.101341e-10, 6.641301e-10, 
    7.181228e-09, 7.718228e-09, 3.180605e-08, 9.611796e-09, -7.489803e-09, 
    7.928946e-09, 1.345862e-08, 4.567056e-09, -1.361485e-09, -9.885071e-11, 
    -9.899736e-09, -3.606999e-11, -6.206591e-12, -1.024333e-08, -8.47018e-10, 
    1.194871e-09, -1.896069e-09, -1.021277e-09, -6.83285e-10, -8.65677e-09, 
    4.038412e-09, -2.353848e-08, -6.064411e-10, 8.172435e-10, 9.381651e-11, 
    4.708056e-10, -1.415685e-09, 8.435563e-10, 1.308592e-10, -2.44782e-12, 
    -5.358913e-11, -8.928851e-09, -1.869192e-08, -2.077722e-08, 
    -1.633389e-09, 7.116796e-11, -1.773515e-09, -1.793154e-09, -1.262754e-08, 
    4.447657e-09, -1.16583e-09, 1.230768e-08, -1.07359e-08, -1.582492e-08, 
    2.139899e-09, 1.402128e-09, 8.100756e-10, -5.541665e-10, 4.659853e-09, 
    1.380673e-09, 1.470823e-10, 1.861267e-11, -2.366363e-09, -3.652168e-10, 
    -5.974528e-10, 3.8699e-10, 8.0028e-10, -1.29603e-10, 1.195778e-08, 
    -6.343782e-09, 3.158107e-09, -2.454527e-09, 1.670628e-10, -6.118568e-10, 
    -1.798924e-09, 7.571089e-09, -1.117769e-09, 7.065637e-11, 5.114877e-09, 
    -1.252886e-09, -1.513345e-08, 9.302426e-11, 4.708653e-09, 3.011849e-10, 
    -4.143317e-11, -1.450502e-09, 3.202061e-11, -1.844986e-09, 1.291873e-10, 
    5.576908e-10, 5.104539e-10, 1.333461e-09, 2.145896e-09, -1.492111e-09, 
    1.215756e-08, 1.650733e-10, 8.154188e-11, -1.210992e-09, -1.293358e-09, 
    -1.117286e-09, 1.42731e-10, 2.271605e-11, 2.827871e-11, -1.495106e-10, 
    -7.979679e-10,
  -6.377832e-11, 2.682839e-09, 3.175501e-09, -7.517826e-10, 2.005862e-09, 
    1.941459e-09, 5.080523e-09, -1.14191e-08, -6.489245e-09, 1.498847e-09, 
    7.366623e-10, -7.456435e-09, 2.131486e-09, -1.97366e-09, -4.475169e-09, 
    -7.387113e-10, -8.708346e-09, 1.484722e-09, -4.087255e-10, 7.947563e-10, 
    -1.163073e-09, 1.534431e-09, 8.328414e-10, 2.013394e-10, -7.203482e-10, 
    6.965564e-09, 6.248371e-09, 4.327913e-08, -1.105403e-08, -4.619721e-09, 
    1.193786e-08, 1.184853e-08, 8.114284e-09, -3.336908e-09, -1.057288e-11, 
    -1.44515e-08, -4.514419e-10, 2.085443e-11, -5.717453e-09, -1.024077e-09, 
    2.162136e-09, -1.202977e-09, -2.049582e-09, -6.474634e-10, -7.824752e-09, 
    2.982119e-09, -2.451424e-08, -6.921042e-10, 6.223388e-10, 8.550671e-11, 
    -9.52646e-10, -2.048751e-09, 1.383665e-09, 2.577622e-10, 2.213767e-11, 
    -3.865352e-12, -1.380528e-08, -2.725494e-08, -9.232329e-09, 
    -5.285816e-09, -1.011387e-09, -6.672565e-10, -1.631037e-09, -1.87218e-08, 
    -1.999871e-09, -1.525478e-09, 1.467524e-08, -1.700832e-08, -1.09633e-08, 
    -1.381463e-08, 7.984511e-10, 8.029133e-11, 2.356046e-09, 5.163201e-09, 
    3.319315e-10, 2.673914e-10, 2.755485e-11, -2.918334e-09, -4.737331e-10, 
    -7.008481e-09, 1.682707e-10, 1.479829e-09, -2.907541e-11, 7.825918e-09, 
    4.445099e-09, 2.207514e-09, 4.993638e-09, 2.484057e-10, -2.176882e-09, 
    -3.922125e-09, 6.07875e-09, -4.686171e-10, 2.45457e-10, 5.256716e-09, 
    2.99616e-09, -2.30199e-08, 2.30068e-10, 3.997741e-09, 1.434046e-09, 
    -9.825953e-11, 1.452634e-10, 1.782823e-10, -2.603413e-09, 1.856488e-10, 
    9.288783e-10, 7.835013e-10, -2.380318e-10, 3.334151e-10, -2.559148e-09, 
    1.655292e-08, 4.866649e-10, 2.773959e-11, -2.442277e-10, -2.489713e-09, 
    -1.398206e-09, 1.466418e-10, 8.682122e-11, -3.368861e-11, -1.278284e-10, 
    -2.335696e-10,
  -5.312017e-10, -1.127887e-09, 1.283809e-09, -1.962803e-09, -4.579306e-10, 
    -4.342837e-10, 4.951062e-10, -1.32593e-09, -1.428475e-08, 3.471428e-10, 
    -1.33133e-09, -1.01478e-08, 5.149445e-09, 2.166757e-09, -5.803429e-09, 
    7.945173e-10, -5.671694e-09, 1.880636e-09, -2.061761e-09, 7.457288e-10, 
    -1.230887e-09, 1.669548e-09, 1.940634e-09, 4.716867e-10, -2.764864e-10, 
    -2.144418e-09, 1.585443e-08, -6.841049e-09, -3.9057e-08, -9.677024e-10, 
    1.528161e-08, 1.045362e-08, 1.339811e-08, -3.538162e-09, -5.027744e-09, 
    -1.689762e-08, -9.967324e-10, 4.641265e-11, 1.212085e-07, -1.103337e-09, 
    4.548031e-09, 4.075105e-10, -3.009234e-09, -5.43765e-10, -2.093202e-09, 
    1.940293e-09, -2.265969e-08, -1.156167e-09, 2.7851e-10, 1.496758e-11, 
    -1.800906e-09, -3.715058e-09, 1.845967e-09, 5.464472e-10, 5.74488e-11, 
    7.426593e-11, -2.439106e-08, -3.56439e-08, 1.728496e-08, -1.249211e-08, 
    -2.48059e-09, 6.856453e-10, -8.341772e-10, -1.788242e-08, -1.671949e-08, 
    -1.770672e-10, 1.703609e-08, -2.10627e-08, -1.58019e-08, -1.811713e-08, 
    -1.65403e-09, 8.130314e-10, 2.519357e-09, 1.910394e-09, -2.433046e-09, 
    4.222329e-10, 6.028245e-11, -3.850985e-09, -6.303523e-10, -6.682853e-09, 
    -9.436292e-10, 4.040589e-09, -2.029594e-10, 5.397339e-09, 6.500272e-09, 
    1.221679e-09, 3.290609e-09, 3.549872e-10, -4.50655e-09, -6.811604e-09, 
    8.4666e-09, 9.848655e-11, 2.447393e-10, 2.775778e-09, 6.010112e-09, 
    -2.904063e-08, -6.957173e-10, 7.770439e-09, 2.440288e-09, -1.368335e-10, 
    -9.737278e-10, 2.04313e-10, -2.700414e-09, 2.833112e-10, 3.89889e-09, 
    1.92955e-09, -7.765948e-10, -5.890001e-09, 1.7763e-09, 1.429811e-08, 
    1.051035e-10, -5.953211e-10, 3.768264e-09, -4.320327e-09, -3.005766e-09, 
    7.339622e-11, 1.646043e-10, -1.112976e-10, -9.434942e-11, 1.648459e-11,
  -1.19087e-10, -3.989044e-09, -1.328203e-09, -1.525848e-09, -1.957631e-09, 
    -1.156991e-09, -3.651849e-09, 6.164612e-09, -1.699709e-08, -7.624351e-09, 
    -7.857977e-09, -1.110254e-08, 3.992739e-09, 1.028803e-08, -3.450907e-09, 
    2.629776e-09, -4.426278e-09, 3.889511e-10, -4.23843e-09, 1.996341e-10, 
    2.672778e-10, 8.192274e-10, 2.822787e-09, 1.068372e-09, 6.412506e-10, 
    6.522214e-10, 2.730604e-08, 2.283286e-09, -4.188513e-08, 9.276619e-09, 
    1.788328e-08, 9.812311e-09, 2.194167e-08, -6.596508e-09, -1.160322e-08, 
    -1.421517e-08, -3.218571e-09, 2.928857e-11, 9.729814e-08, -1.43221e-09, 
    9.682855e-09, 2.957961e-09, -3.777473e-09, -1.116651e-09, -2.413401e-09, 
    3.462901e-10, -2.906216e-08, -2.950955e-09, -1.664603e-09, -6.671286e-11, 
    -8.58762e-10, -6.386188e-09, 2.55767e-09, 1.076933e-09, 2.181764e-10, 
    1.157048e-10, -2.731912e-08, -4.224256e-08, 3.544471e-08, -2.156106e-08, 
    -5.155073e-09, 9.625296e-10, -2.045226e-10, -1.152282e-08, -2.648267e-08, 
    -1.666649e-10, 2.095118e-08, -2.223595e-08, -1.627882e-08, -7.648737e-09, 
    -2.441277e-08, 1.260071e-08, -1.555622e-08, 8.845404e-10, -3.865608e-09, 
    7.280505e-10, 1.154348e-10, -4.636249e-09, -8.16577e-10, -3.783043e-09, 
    -2.68895e-09, 8.296372e-09, -7.54028e-10, -1.026365e-09, 9.435098e-09, 
    1.223384e-09, -1.983835e-11, 8.117809e-10, -7.733818e-09, -1.010068e-08, 
    1.039928e-08, 1.052239e-09, -2.471552e-10, -6.182646e-09, 9.918779e-09, 
    -4.115007e-08, -1.948127e-09, 1.549239e-08, 3.231492e-09, -2.575575e-10, 
    -1.591332e-09, -1.329852e-10, -3.26261e-09, 4.301555e-10, 8.38395e-09, 
    8.323752e-09, 3.490186e-11, -1.475007e-08, 1.230819e-08, 7.634924e-09, 
    -1.256012e-09, -1.790283e-09, 8.050563e-09, -3.686182e-09, -1.330534e-08, 
    4.638992e-11, 3.755645e-10, -1.299387e-10, -6.953726e-11, -1.979856e-10,
  4.366143e-10, -8.175789e-10, -1.87265e-09, -4.16378e-10, -1.821263e-09, 
    -1.362366e-09, -2.633612e-09, 4.508991e-09, -6.343896e-09, -2.993988e-08, 
    -1.537734e-08, -1.106963e-08, -1.145906e-09, 8.704092e-09, 7.061431e-09, 
    1.149653e-09, -5.36707e-09, -2.651205e-09, -5.963898e-09, -1.038302e-09, 
    1.838544e-09, 2.139586e-10, 1.970363e-09, 2.058641e-09, -2.90413e-10, 
    2.830802e-09, 2.445091e-08, 1.316005e-08, -5.093813e-08, 1.339009e-08, 
    1.996983e-08, 1.205586e-08, 2.839158e-08, -1.042741e-08, -3.259458e-09, 
    -1.142394e-08, -5.391769e-09, 4.174439e-11, 1.776164e-08, 2.003833e-09, 
    2.538023e-08, 4.542187e-09, -4.455288e-09, -4.008706e-09, -8.226948e-09, 
    2.131173e-09, -4.539996e-08, -2.736797e-09, -6.502091e-09, -1.166285e-10, 
    -2.645983e-09, -9.857388e-09, 4.079777e-09, 1.980993e-09, 5.536123e-10, 
    1.122089e-10, -3.7169e-08, -4.864627e-08, 9.761027e-09, -2.91073e-08, 
    -3.048626e-09, -1.500666e-10, -9.111432e-10, -3.16802e-09, -2.759757e-08, 
    -1.817e-09, 2.936707e-08, -2.003446e-08, -1.853954e-08, -1.705934e-08, 
    -6.948909e-08, 4.072973e-08, -2.699051e-08, -3.068067e-09, -3.271623e-09, 
    1.179615e-09, 5.665157e-11, -4.942621e-09, -1.0189e-09, -4.246203e-11, 
    -5.391882e-09, 1.22232e-08, -1.358245e-09, 1.0902e-09, 5.725951e-09, 
    1.410683e-09, -3.061757e-09, 1.926878e-09, -1.289393e-08, -1.566499e-08, 
    8.582958e-09, 2.850902e-09, -1.001581e-09, -1.26553e-08, 1.299333e-08, 
    -7.012299e-08, -5.008166e-09, 1.483227e-08, 5.43082e-09, -5.011657e-10, 
    -1.248168e-09, -8.15394e-10, -4.053526e-09, 6.834604e-10, 1.166728e-08, 
    7.38811e-09, -3.667537e-10, -1.333461e-08, 1.731809e-08, 1.644992e-09, 
    -6.86498e-10, -4.009223e-09, 9.678104e-09, -8.382699e-10, -2.832456e-08, 
    8.802772e-11, 7.037571e-10, -1.139089e-10, -7.641532e-11, -1.955982e-10,
  2.912657e-10, 8.219558e-11, -7.368612e-10, -2.981437e-10, -5.441052e-10, 
    -6.75243e-10, 2.219451e-09, -3.287937e-09, 3.024923e-09, -1.794052e-08, 
    -1.973683e-08, -1.037728e-08, -7.729909e-09, 3.537764e-09, 1.677415e-08, 
    -1.834479e-09, -5.289553e-09, -4.21727e-09, -4.125582e-09, -1.988099e-09, 
    1.078206e-09, 3.002697e-09, -3.553851e-10, 3.352e-09, -9.831638e-10, 
    2.708703e-09, 4.982269e-08, 3.553646e-08, -5.279213e-08, -1.322519e-08, 
    2.20756e-08, 1.660226e-08, 2.759225e-08, -1.684708e-08, 7.139477e-09, 
    -6.891412e-09, -7.77556e-09, 6.617995e-11, -4.202434e-10, 5.76299e-09, 
    3.360189e-08, 3.62428e-09, -6.04598e-09, -2.352845e-09, 1.617423e-09, 
    2.498041e-09, -4.964483e-08, -2.698357e-09, -1.258742e-08, -2.181899e-10, 
    -1.956636e-09, -1.261151e-08, 6.081183e-09, 3.42709e-09, 1.205107e-09, 
    6.08793e-11, -4.887852e-08, -5.654207e-08, -5.830249e-08, -4.535567e-08, 
    2.023114e-09, -2.065462e-09, -1.067122e-09, 1.040055e-08, -2.91756e-08, 
    -1.973206e-09, 3.080601e-08, -1.715574e-08, -3.329887e-08, -2.110482e-08, 
    -5.827496e-08, 5.107819e-08, -2.223823e-08, -3.024468e-09, -3.275073e-09, 
    1.481055e-09, 9.338663e-11, -4.324704e-09, -1.289821e-09, 8.851089e-10, 
    -1.094475e-08, 1.83196e-08, -1.702631e-09, 8.650431e-10, 5.120455e-10, 
    2.107413e-09, -9.980454e-09, 4.153947e-09, -1.556952e-08, -2.319129e-08, 
    4.461356e-09, 6.000641e-09, -1.998401e-09, -1.395232e-08, 2.031538e-08, 
    -1.199112e-07, -2.829564e-09, -8.944994e-09, 8.268614e-09, -1.003582e-09, 
    -3.901164e-10, -4.633769e-10, -5.51071e-09, 1.053447e-09, 3.527646e-09, 
    1.057913e-09, -9.715166e-09, 3.314256e-09, 1.160566e-08, -1.33582e-10, 
    -2.00032e-10, -4.862045e-09, 1.28756e-09, 7.895892e-09, -6.76431e-09, 
    1.38516e-10, 1.137018e-09, -1.172591e-10, -1.014939e-10, -3.472564e-10,
  -2.761453e-10, 5.200604e-10, -3.897185e-10, -2.166985e-09, -2.39686e-09, 
    -2.683237e-09, 4.325216e-09, -8.828863e-09, 1.198936e-08, -6.22606e-10, 
    -4.726701e-09, -1.888111e-09, -3.707271e-09, -1.048079e-09, 2.087808e-08, 
    -1.657764e-09, -6.160712e-09, -5.539192e-09, 4.741452e-10, -3.399975e-09, 
    -5.877098e-09, 5.740162e-09, 6.513346e-09, 1.383285e-09, -1.135334e-09, 
    9.587779e-10, -1.190227e-08, 3.694635e-08, -3.584978e-08, -2.19448e-08, 
    2.192047e-08, 1.784281e-08, 2.538343e-08, -2.302306e-08, 8.755705e-09, 
    -1.113e-08, -1.262092e-08, 1.590763e-10, 1.418715e-08, 9.940846e-09, 
    1.791675e-08, 1.40119e-10, -8.896251e-09, 1.119054e-08, 7.709843e-09, 
    -4.743811e-09, -5.184071e-08, -1.39228e-09, -1.697847e-08, -3.414904e-10, 
    5.298375e-10, -8.380823e-09, 7.439303e-09, 5.517324e-09, 2.342593e-09, 
    7.503331e-12, -5.045905e-08, -6.583178e-08, -9.351673e-08, -7.802754e-08, 
    -2.232412e-09, -6.365326e-09, -1.725482e-09, 2.600876e-08, -3.239747e-08, 
    5.740617e-10, 3.217497e-08, -1.163346e-08, -5.689299e-08, -2.538604e-08, 
    -2.21707e-08, 4.268333e-08, -2.708634e-08, -2.958132e-09, -6.257642e-09, 
    1.988099e-09, 2.992451e-10, -3.407308e-09, -1.301031e-09, 9.934524e-10, 
    -2.014252e-08, 3.019591e-08, -1.567997e-09, 1.155342e-09, -4.79281e-09, 
    1.867022e-09, -1.776016e-08, 7.005667e-09, -1.771923e-08, -3.212114e-08, 
    7.858034e-10, 9.473695e-09, -2.90909e-09, 7.277876e-10, 3.21624e-08, 
    -1.697409e-07, 1.217769e-08, -2.674221e-08, 8.970687e-09, -1.988519e-09, 
    1.892886e-10, 4.591527e-10, -7.869435e-09, 1.253959e-09, 1.200306e-09, 
    -3.209436e-09, -3.639229e-09, 1.517088e-08, 7.044093e-09, -3.244622e-10, 
    -3.678338e-10, -3.325056e-09, -2.74872e-09, 6.672792e-09, 6.712071e-09, 
    1.370722e-10, 1.320025e-09, -1.222915e-10, -9.205436e-11, -1.428759e-09,
  -3.386731e-10, -2.908109e-10, 2.571028e-10, -3.589946e-09, -4.035599e-09, 
    -5.630568e-09, -7.109975e-10, -9.753592e-09, 1.011114e-08, 1.306006e-08, 
    8.043855e-09, 4.071296e-09, -2.196998e-10, -4.204708e-10, 1.417794e-08, 
    1.218906e-08, -8.966805e-09, -6.662276e-09, 6.692488e-09, -8.890424e-09, 
    -2.061546e-08, -2.825266e-08, -1.960979e-08, -6.718494e-09, 
    -2.936531e-10, 2.763159e-10, -2.159055e-08, -5.247443e-09, -1.489639e-09, 
    -2.835446e-08, 2.441755e-08, 1.662147e-08, 3.542141e-08, -3.035973e-08, 
    4.068681e-09, -2.273805e-08, -1.579643e-08, 2.193943e-10, -2.290847e-09, 
    1.413801e-08, 3.527589e-10, -4.565607e-09, -1.073568e-08, 1.36112e-08, 
    3.978602e-08, -2.219713e-08, -6.375447e-08, 3.055703e-09, -1.921597e-08, 
    -4.779963e-10, 5.072003e-09, 5.399329e-09, 6.165755e-09, 8.840743e-09, 
    3.300752e-09, -1.05274e-10, -6.316964e-08, -7.671115e-08, -8.787052e-08, 
    -5.012387e-08, -1.984063e-09, -4.716753e-09, 8.662937e-11, 3.346442e-08, 
    -2.964973e-08, 7.055519e-09, 4.067169e-08, -1.479691e-09, -7.284586e-08, 
    -2.433586e-08, -4.832344e-08, 2.209123e-08, -3.725552e-08, -2.046704e-09, 
    -2.091962e-08, 2.433126e-09, 2.520295e-10, -2.483375e-09, -1.220053e-09, 
    8.328698e-10, -2.927547e-08, 4.093538e-08, -9.646897e-10, 1.691376e-09, 
    -2.658965e-09, -1.545573e-09, -2.231718e-08, 7.0238e-09, -1.922434e-08, 
    -4.237648e-08, -2.075694e-09, 1.532329e-08, -3.118174e-09, 5.303193e-09, 
    1.648004e-08, -1.629633e-07, 3.954898e-08, 1.556731e-08, 9.473752e-09, 
    -3.811488e-09, 5.109086e-10, 7.985292e-10, -1.057629e-08, 3.24146e-10, 
    -1.517435e-09, 5.95719e-10, 5.067079e-09, 1.394773e-08, 2.907143e-09, 
    -1.029264e-09, -2.180798e-09, -4.702656e-10, -1.42569e-09, 2.093543e-09, 
    1.494732e-08, -9.464429e-12, 1.440497e-09, -1.073559e-10, -7.261747e-12, 
    -1.891976e-09,
  -1.559215e-10, -3.46347e-10, 1.894307e-09, -1.604519e-09, -3.98353e-09, 
    -5.305594e-09, -5.839581e-09, -7.789765e-09, -3.4766e-09, 1.50697e-08, 
    1.290215e-08, 2.311992e-09, 1.038529e-10, -1.154092e-09, -1.751289e-09, 
    2.800091e-08, -1.502175e-08, -8.03243e-09, 1.347878e-08, -1.88241e-08, 
    -3.139218e-08, -5.13532e-08, -5.000624e-08, -1.456857e-08, 7.362928e-10, 
    1.170463e-09, -1.570584e-10, -1.773952e-08, 1.635436e-08, -4.399539e-08, 
    3.590202e-08, 1.499103e-08, 6.10857e-08, -3.824738e-08, 1.395506e-10, 
    -4.682516e-08, -1.776796e-08, 2.036415e-10, -2.239693e-08, 1.784449e-08, 
    -1.402158e-08, -2.939885e-09, -1.088193e-08, 8.640816e-09, 6.160116e-08, 
    -7.420243e-08, -7.701294e-08, 5.874966e-09, -2.25241e-08, -6.277787e-10, 
    1.304166e-08, -1.889532e-09, 9.79594e-10, 1.153879e-08, 2.553182e-09, 
    -1.836611e-10, -6.654142e-08, -8.869569e-08, -8.025509e-08, 
    -2.062333e-08, 3.786397e-09, -1.35384e-09, 2.822674e-09, 2.219118e-08, 
    -2.733863e-08, 9.950952e-09, 4.499378e-08, 1.018572e-08, -6.398062e-08, 
    -1.154996e-08, -7.693353e-08, 6.835421e-10, -5.788235e-08, 2.747299e-09, 
    -5.577709e-08, -1.311776e-09, -6.698428e-10, -1.895444e-09, 
    -1.055645e-09, 3.12923e-10, -3.500224e-08, 3.700929e-08, -1.465992e-10, 
    1.33565e-09, -1.10191e-09, -5.193044e-09, -1.031918e-08, 4.987498e-09, 
    -2.007903e-08, -5.127026e-08, -6.899711e-09, 1.263126e-08, -3.179707e-09, 
    2.997751e-08, 2.013564e-09, -1.035731e-07, 5.786977e-08, 3.291115e-08, 
    5.649724e-09, -6.04665e-09, -4.015988e-10, -9.303086e-09, 1.35622e-09, 
    -1.476153e-09, -5.25705e-09, 3.823345e-09, -4.198398e-09, 5.680874e-09, 
    6.511414e-10, -2.69182e-09, -4.74364e-09, 2.689262e-10, 1.402327e-10, 
    -8.206996e-09, 5.908134e-09, 2.671641e-11, 1.424368e-09, -2.552767e-10, 
    2.080469e-11, 4.999379e-10,
  6.548362e-11, -1.11072e-10, 3.186074e-09, 4.61057e-09, -4.215053e-09, 
    -4.36512e-09, -5.060201e-09, -4.849767e-09, -1.493459e-08, 5.017682e-09, 
    5.831225e-09, -1.40858e-10, -1.762146e-10, -1.558305e-09, -1.158469e-09, 
    4.306112e-08, -1.970909e-08, -1.034829e-08, 2.088787e-08, -3.27143e-08, 
    -2.67288e-08, -3.801949e-08, -4.45383e-08, -1.237322e-08, -9.920313e-10, 
    3.082846e-09, -2.583351e-08, -1.016588e-08, 4.438448e-09, -7.819688e-08, 
    2.812283e-08, 2.641957e-08, 8.058953e-08, -3.272771e-08, 4.832827e-09, 
    -9.901123e-08, -1.844168e-08, 5.169909e-11, -1.837373e-08, 2.164178e-08, 
    -3.409421e-08, 4.322828e-09, -1.147484e-08, 3.049632e-10, 3.42103e-08, 
    -1.466597e-07, -8.642508e-08, 1.198831e-08, -2.057038e-08, -2.115947e-09, 
    1.807435e-08, -1.75105e-08, -5.817026e-09, 1.408703e-08, -1.601563e-11, 
    -3.075229e-10, -6.706443e-08, -9.395641e-08, -1.057273e-07, 
    -1.321409e-08, 8.776055e-09, 2.042157e-09, 1.682565e-09, 3.142274e-08, 
    -6.455745e-08, 7.169433e-09, 2.730928e-08, 1.864885e-08, -3.043363e-08, 
    -3.166747e-09, -8.650522e-08, -8.912366e-09, -3.981904e-08, 4.347726e-09, 
    -7.165016e-08, -7.796984e-09, -1.327635e-09, -2.650523e-09, 
    -1.989724e-09, 5.734364e-10, -3.898953e-08, 1.52892e-08, 1.153353e-10, 
    -7.25322e-10, -8.038796e-10, 1.049898e-09, -1.73543e-09, 3.35433e-09, 
    -3.043664e-08, -5.887131e-08, -9.635414e-09, 4.67826e-09, -1.723635e-09, 
    9.855086e-08, -3.145044e-08, -6.5279e-08, 6.94602e-08, 1.983608e-09, 
    1.002491e-09, -7.586868e-09, -2.835577e-09, -3.636806e-08, 1.20896e-08, 
    -2.658957e-09, -2.144134e-09, 7.06757e-09, -8.357802e-09, 6.476512e-09, 
    1.267608e-09, -3.349669e-09, -5.733114e-09, 2.127081e-10, 1.319449e-09, 
    -2.02499e-08, -9.879386e-11, -6.631353e-11, 1.625708e-09, -2.407745e-10, 
    1.332126e-10, 3.105924e-09,
  6.417054e-10, -3.359446e-11, 2.144645e-09, 1.55573e-08, -3.308571e-09, 
    -4.034462e-09, -4.857554e-09, -4.667413e-10, -1.104496e-08, -1.02761e-08, 
    -2.285674e-10, -3.666969e-10, 1.249703e-09, -5.030245e-09, -2.35417e-09, 
    5.380384e-08, -1.586279e-08, -1.71176e-08, 3.08914e-08, -4.634802e-08, 
    6.620724e-09, -2.112625e-08, -1.57948e-08, -2.472808e-08, -9.571806e-09, 
    4.974197e-09, -2.527423e-08, -2.226727e-09, -1.569055e-08, -9.38698e-08, 
    4.980762e-08, 4.99486e-08, 7.971033e-08, -1.521067e-08, 4.619665e-10, 
    -1.478433e-07, -1.847097e-08, -4.184244e-10, -8.468589e-09, 9.955112e-09, 
    -5.993135e-08, 2.918625e-09, -9.554924e-09, -1.358004e-08, 3.16773e-08, 
    -1.268984e-07, -8.709191e-08, 1.331347e-08, -1.34021e-08, 1.03654e-09, 
    2.048455e-08, -1.056122e-08, -1.110436e-08, 1.689749e-08, -2.035833e-09, 
    -3.981881e-10, -9.080389e-08, -8.124455e-08, -1.79398e-07, -1.488776e-08, 
    6.427797e-09, 1.588603e-09, -9.941914e-11, 5.834255e-08, -8.712536e-08, 
    2.087705e-08, -1.382779e-08, 2.58745e-08, -1.744894e-08, 2.122221e-08, 
    -1.686417e-07, 1.761578e-10, -1.118775e-08, 1.860883e-09, -5.130939e-08, 
    -1.288566e-08, -1.62197e-09, -7.36614e-09, -2.345317e-09, -2.966658e-10, 
    -4.662706e-08, -1.083384e-08, -9.032419e-11, -2.24594e-09, -3.261505e-09, 
    -6.148468e-09, 7.877532e-09, 1.948194e-09, -4.643997e-08, -6.778828e-08, 
    -6.410062e-09, 9.928078e-09, 6.642153e-10, 1.610546e-07, -2.168377e-08, 
    -3.625621e-08, 8.468099e-08, 2.720583e-09, -7.23702e-09, -8.074823e-09, 
    -2.987741e-08, -5.58951e-08, 1.735506e-08, -4.211181e-09, -1.076899e-09, 
    2.326846e-08, -5.084701e-09, 1.5696e-08, 4.918377e-09, -3.428227e-10, 
    -5.720437e-09, 6.404548e-10, 1.558078e-10, -2.234577e-08, -4.985168e-11, 
    2.649699e-10, 1.520903e-09, -3.614957e-10, 2.692673e-10, 6.89937e-09,
  1.56939e-09, -9.589485e-11, 1.027104e-09, 1.102904e-08, -2.957563e-10, 
    -3.730577e-09, -4.959759e-09, -1.247656e-09, 2.153854e-09, -1.073619e-08, 
    -9.76371e-09, -2.370541e-09, 3.223022e-11, -1.583334e-08, 1.064052e-09, 
    6.052552e-08, -5.253231e-09, -2.098818e-08, 4.363618e-08, -5.806231e-08, 
    5.377075e-08, -2.283019e-08, -3.380649e-09, -1.398433e-08, -8.957329e-09, 
    1.367596e-09, 1.01444e-07, 6.02671e-09, -1.317147e-08, -7.653802e-08, 
    2.357461e-08, 2.656128e-08, 3.72201e-08, 1.490099e-08, 7.975132e-11, 
    -1.525936e-07, -2.49605e-08, -1.097661e-09, -1.68655e-08, 2.468093e-08, 
    -8.462727e-08, 2.561933e-10, -9.364129e-09, -3.523732e-08, 4.730492e-08, 
    -4.353598e-08, -6.719108e-08, 3.322043e-09, -1.496379e-08, 7.070447e-09, 
    2.088184e-08, -1.127279e-08, -1.020492e-08, 2.081632e-08, -4.863261e-09, 
    -3.645368e-10, -7.593093e-08, -4.667593e-08, -2.406346e-07, 
    -2.189721e-08, 3.113371e-09, 7.395329e-11, -6.797904e-10, 9.16673e-08, 
    -8.906191e-08, 2.186977e-08, -3.991903e-08, 4.334396e-08, -3.815529e-08, 
    4.695124e-08, -1.929631e-07, 2.830865e-08, 4.360743e-09, 8.93408e-10, 
    -1.818766e-08, -1.593668e-08, -1.358188e-09, -1.341434e-08, 
    -3.153846e-09, -2.776972e-09, -5.320106e-08, -2.676352e-08, 1.995204e-11, 
    -3.440334e-09, -1.716984e-08, 5.375512e-09, 9.913663e-09, 1.659657e-09, 
    -6.738597e-08, -9.028668e-08, -8.35314e-10, 1.00894e-08, 3.146425e-09, 
    2.054091e-07, -2.658254e-08, -1.202147e-08, 1.108177e-07, -3.66685e-08, 
    -1.899053e-08, -8.70674e-09, -4.108364e-08, -5.134837e-08, 2.137514e-08, 
    -5.702375e-09, 1.400502e-08, 2.323037e-08, 2.807212e-09, 2.51726e-08, 
    8.966083e-09, 2.100649e-09, -7.433414e-10, 1.434216e-09, -3.245816e-09, 
    -1.928976e-08, 3.084835e-09, 3.453351e-10, 1.293742e-09, -2.720313e-10, 
    3.725162e-10, 1.194468e-08,
  1.160515e-09, -2.694378e-11, 1.008175e-09, 3.561695e-09, 2.324896e-10, 
    -2.430511e-09, -4.456751e-09, -3.894229e-09, -6.399091e-09, 
    -4.981075e-09, -6.545974e-09, -4.455728e-09, 9.839596e-10, -9.860628e-09, 
    3.485411e-09, 5.702948e-08, 1.821672e-09, -2.543186e-08, 5.766732e-08, 
    -7.199446e-08, 8.415714e-08, -4.070307e-08, -9.018322e-09, 5.263701e-09, 
    7.929657e-10, -1.495209e-09, 3.89167e-07, 4.978347e-10, 3.708578e-09, 
    -6.191488e-08, -4.19177e-08, -2.618322e-09, -2.969455e-08, 1.326623e-08, 
    2.109459e-09, -1.18508e-07, -3.939775e-08, -1.67995e-09, -2.904426e-08, 
    3.045675e-08, -9.44955e-08, 4.968115e-11, 6.193403e-09, -5.047877e-08, 
    4.523781e-08, 2.21462e-08, -3.862203e-08, -2.187176e-08, -1.659382e-08, 
    1.298474e-08, 1.986854e-08, -1.425178e-09, -7.787571e-09, 2.612023e-08, 
    -7.215115e-09, -1.163585e-10, -6.552239e-08, -4.391165e-09, 
    -2.848347e-07, -1.958189e-08, 3.316472e-09, -4.963567e-10, -6.898517e-10, 
    1.064186e-07, -2.86384e-08, -7.368953e-09, -3.769435e-08, 2.496608e-07, 
    -8.001143e-08, 6.670462e-09, -2.138567e-07, 2.090076e-08, 7.697508e-09, 
    -1.750209e-09, 5.330162e-09, -9.023552e-09, -1.317702e-09, -1.661653e-08, 
    -3.750301e-09, -7.192614e-08, -8.906164e-08, -4.145608e-08, 2.659533e-09, 
    -3.485184e-09, -1.955527e-08, -5.116021e-08, -6.818823e-09, 
    -1.190642e-09, -9.336418e-08, -1.262521e-07, 5.216634e-09, -3.090713e-09, 
    3.791428e-09, 2.143654e-07, -6.383675e-08, 1.206655e-08, 1.516322e-07, 
    -7.239919e-09, -3.282264e-08, -1.02915e-08, -1.805915e-09, -2.711989e-08, 
    2.716744e-08, -7.709154e-09, 3.817649e-08, 3.136654e-08, 2.056584e-08, 
    2.157435e-08, 1.258547e-08, 1.595367e-09, 9.653377e-09, 4.772573e-10, 
    -6.736514e-09, -1.620356e-08, 2.858656e-09, 2.291699e-10, 7.229772e-10, 
    -4.238991e-10, 4.239027e-10, 9.08733e-09,
  -6.819903e-09, -3.029754e-11, 8.894006e-09, 1.611619e-08, 4.428841e-09, 
    2.677837e-09, -9.00684e-10, -2.269473e-09, -1.507232e-08, -7.735537e-09, 
    -4.265246e-09, -1.249816e-09, 1.687056e-09, -8.009181e-09, 1.402685e-08, 
    3.568431e-08, 2.053295e-08, -3.058551e-08, 7.298549e-08, -8.910314e-08, 
    8.356659e-08, -5.460203e-08, -1.482618e-08, 6.904031e-09, 4.142123e-09, 
    3.577156e-10, 1.94651e-07, 1.345524e-08, 3.617487e-08, -5.842986e-08, 
    -4.448117e-08, -9.896269e-09, -5.652345e-08, 2.71138e-08, 5.082768e-09, 
    -5.287626e-08, -6.278186e-08, -1.956153e-09, -5.623684e-08, 5.931433e-08, 
    -7.047503e-08, 3.115588e-10, 1.64124e-08, -5.533681e-08, 3.066629e-08, 
    5.258454e-08, -2.131361e-08, -3.192355e-08, -7.509799e-09, 1.337376e-08, 
    1.813527e-08, -3.615963e-08, -9.622783e-09, 3.401959e-08, -1.050162e-08, 
    -1.215824e-09, -7.438149e-08, 1.053463e-08, -3.511863e-07, -2.132472e-08, 
    6.604694e-09, -6.891128e-10, -3.017817e-10, 1.281961e-07, 4.513419e-08, 
    2.025655e-08, -6.503984e-08, 2.851451e-07, -7.350076e-08, 2.275726e-09, 
    -2.396103e-07, -3.035854e-08, -2.222731e-08, 2.814943e-09, 2.102337e-08, 
    -6.203948e-09, -2.287791e-09, -1.772128e-08, -4.275546e-09, 
    -1.932851e-07, -1.358918e-07, -5.16644e-08, 7.442736e-09, 4.379956e-09, 
    -1.685123e-09, -1.131164e-07, -4.535451e-08, -1.115211e-09, 
    -1.239333e-07, -1.703011e-07, 3.541516e-09, -1.900952e-08, 3.58736e-09, 
    2.070305e-07, -6.66891e-08, 4.724492e-08, 1.640041e-07, 1.284667e-08, 
    -4.530301e-08, -1.1231e-08, 5.465648e-08, 2.966203e-09, 1.61094e-08, 
    -9.30423e-09, 5.518984e-09, 5.114072e-08, 7.131973e-09, 2.587313e-08, 
    1.614654e-08, -3.854552e-10, 1.314157e-08, -7.244694e-10, -9.762573e-09, 
    -1.557879e-08, 3.621437e-09, 8.444431e-10, 2.99849e-10, -1.21106e-09, 
    4.849596e-10, 6.079006e-09,
  -3.307628e-08, 2.657998e-10, 1.955016e-08, 2.810543e-08, 7.786525e-09, 
    8.331881e-09, -1.968942e-09, -1.297281e-09, -1.148294e-08, 3.685386e-09, 
    -3.62661e-10, 6.65068e-10, 9.370069e-10, 2.623551e-09, 2.358661e-09, 
    2.630918e-08, 2.061397e-08, -3.259447e-08, 8.444735e-08, -9.316705e-08, 
    5.077743e-08, -3.442233e-08, -1.502201e-08, 1.925059e-09, 5.527909e-09, 
    1.369244e-09, 1.316369e-08, 3.237653e-08, 2.215052e-08, -4.424612e-08, 
    5.30315e-09, 9.903829e-09, -3.731282e-08, 5.356765e-08, 5.493916e-09, 
    -2.315915e-09, -9.135366e-08, -3.057636e-09, -8.898166e-08, 9.081355e-08, 
    -1.447554e-08, -1.203603e-09, -1.299617e-08, -5.439522e-08, 1.881438e-08, 
    5.499021e-08, -1.639961e-08, -3.705097e-08, -1.372723e-08, 8.673034e-09, 
    1.625958e-08, -9.055032e-08, -1.57857e-08, 4.347999e-08, -1.473901e-08, 
    2.663683e-10, -1.038868e-07, 1.559864e-08, -3.639661e-07, -2.989222e-08, 
    6.80177e-09, -8.81073e-10, -2.188642e-08, 1.54471e-07, 1.109746e-07, 
    1.100489e-08, -9.893859e-08, 8.405902e-08, -7.069104e-08, 2.141292e-09, 
    -1.831919e-07, -4.365245e-08, -7.43936e-08, 8.527422e-09, 1.868304e-08, 
    -3.253774e-08, -2.759464e-09, -1.553437e-08, -4.008538e-09, 
    -6.355219e-08, -1.817668e-07, -5.697941e-08, 5.337029e-09, 1.09676e-08, 
    8.774464e-09, 1.864453e-08, 3.761601e-07, 2.676188e-10, -1.580849e-07, 
    -2.128883e-07, 7.939889e-10, -2.929796e-08, 5.730612e-09, 1.881877e-07, 
    -3.910748e-08, 1.058483e-07, 1.163125e-07, 2.539298e-08, -5.957236e-08, 
    -1.139633e-08, 1.610852e-08, 2.296822e-08, -3.711833e-09, -1.052994e-08, 
    4.915478e-09, 1.020987e-08, -5.641482e-09, 2.89906e-08, 3.451078e-08, 
    -4.96334e-09, 4.6781e-09, 4.203912e-09, -9.412474e-09, -1.48774e-08, 
    5.639663e-09, 1.916862e-09, 6.842527e-10, -1.303267e-09, 5.719727e-10, 
    -1.399633e-08,
  -4.211552e-08, 1.871626e-09, 1.730882e-08, 2.801994e-08, 8.644406e-09, 
    8.850748e-09, -1.548528e-09, 1.619355e-09, -1.170213e-08, -7.140329e-09, 
    7.008339e-09, 1.349918e-09, 5.494371e-09, -7.25322e-09, 1.587705e-08, 
    2.340706e-08, 2.13839e-08, -3.321645e-08, 9.098618e-08, -5.925642e-08, 
    7.780955e-09, 6.396931e-09, -1.093929e-08, 1.440412e-10, 2.796696e-10, 
    2.110119e-08, -6.342475e-09, 1.122612e-08, 4.006176e-08, -1.870364e-08, 
    9.290147e-09, 2.392949e-08, -1.904505e-08, 1.657872e-08, -3.164928e-09, 
    1.237083e-08, -1.040449e-07, -3.306312e-09, -1.045297e-07, 1.191558e-07, 
    5.040283e-08, -2.947331e-09, -6.136105e-09, -5.294934e-08, 1.686203e-08, 
    4.484275e-08, -2.597523e-08, -4.039674e-08, -2.03311e-08, 3.11632e-09, 
    1.463921e-08, -1.457593e-07, -3.319056e-08, 5.16289e-08, -2.212678e-08, 
    9.225687e-11, -1.356254e-07, 1.120435e-07, -3.790393e-07, -3.528625e-08, 
    3.499849e-09, 7.541189e-09, -1.200622e-07, 1.939925e-07, 9.691502e-08, 
    8.417589e-08, -1.02178e-07, -1.393414e-08, -6.693199e-08, -2.265892e-09, 
    -6.952337e-08, -1.003241e-08, -9.411588e-08, 1.523858e-09, 1.069334e-08, 
    -2.660522e-08, -3.894087e-09, -6.856737e-09, -3.569715e-09, 
    -5.627498e-11, -2.275309e-07, -5.950574e-08, -2.991175e-08, 7.661583e-09, 
    -1.360831e-09, -2.948411e-08, 3.755451e-08, 2.127422e-09, -1.906246e-07, 
    -2.631811e-07, -1.108322e-08, -4.105277e-08, 9.577974e-09, 1.751406e-07, 
    -2.167496e-08, 1.895994e-07, 6.634673e-08, 3.68658e-08, -7.287804e-08, 
    -1.094863e-08, -4.965023e-08, 1.750123e-08, 1.178819e-09, -1.089359e-08, 
    1.626654e-08, -3.0352e-08, 5.125344e-09, 6.152163e-09, 5.369566e-08, 
    -1.457192e-08, 6.889422e-11, 1.277874e-08, 2.839897e-09, -1.2123e-08, 
    5.438437e-09, 2.553133e-09, -6.266703e-10, -1.467107e-09, 6.645919e-10, 
    -4.82944e-08,
  -1.881784e-08, 6.451444e-09, 5.853678e-09, 1.527889e-08, 3.686807e-09, 
    2.38191e-09, -1.035744e-09, 3.634739e-09, -2.097573e-08, -7.574209e-08, 
    1.345086e-09, 1.389196e-09, -2.12728e-08, -3.153383e-08, 3.594363e-08, 
    1.805109e-08, 4.462144e-08, -4.156021e-08, 8.800518e-08, -1.507584e-08, 
    -3.49151e-08, 2.06532e-08, -9.971416e-09, 6.927507e-10, -1.543918e-08, 
    4.801922e-08, -1.375594e-08, 1.415168e-08, 4.82782e-08, -9.683106e-09, 
    4.490232e-09, 3.500685e-08, 4.619665e-10, -6.25181e-09, 2.649529e-09, 
    1.322263e-08, -8.246557e-08, -3.672127e-09, -1.099957e-07, 1.389564e-07, 
    9.425067e-08, -1.336804e-08, -8.954572e-08, -5.430294e-08, 1.041695e-08, 
    2.623625e-08, -4.90075e-08, -4.012844e-08, -2.723105e-08, -4.37602e-10, 
    1.349737e-08, -2.363558e-07, -5.038825e-08, 6.146946e-08, -2.78937e-08, 
    9.083578e-11, -1.424868e-07, -1.088691e-07, -3.87732e-07, -1.982703e-08, 
    2.94159e-09, 2.166831e-08, -2.081355e-07, 2.058909e-07, 7.44048e-08, 
    4.825716e-08, -8.177341e-08, -3.401794e-09, -5.008593e-08, -6.501693e-09, 
    4.235943e-08, 1.84105e-08, -1.15786e-07, -8.359109e-09, 9.928487e-09, 
    -1.750578e-08, -6.925333e-09, -2.784617e-09, -2.730417e-10, 
    -1.883546e-08, -2.570287e-07, -6.99717e-08, -8.345415e-08, -8.957528e-08, 
    -2.858826e-09, -5.720045e-08, -5.766316e-08, 2.399872e-09, -2.166195e-07, 
    -3.122854e-07, 7.095139e-09, -5.037387e-08, 1.133057e-08, 1.814679e-07, 
    -2.07346e-08, 2.652481e-07, 3.219401e-08, 9.134226e-09, -8.43367e-08, 
    -1.343489e-08, -6.525568e-09, -9.23837e-09, -3.856208e-09, -1.053126e-08, 
    1.098903e-08, -2.097846e-08, 5.810756e-08, -1.089558e-08, 5.169869e-08, 
    -2.137784e-08, -6.697462e-09, 1.30421e-08, 2.176154e-08, -9.634107e-09, 
    1.126466e-09, 2.907473e-09, -1.597328e-09, -1.233886e-09, 8.354704e-10, 
    -3.832673e-08,
  1.790227e-09, 2.298202e-08, -9.84744e-09, -2.148454e-09, 8.227289e-09, 
    -7.147037e-09, 2.47735e-09, 4.852723e-09, -2.768888e-08, -9.600069e-08, 
    -6.638425e-08, -1.700244e-08, -1.042645e-08, -4.560502e-08, 1.39413e-08, 
    1.486348e-08, 8.121489e-08, -4.27213e-08, 5.377632e-08, 2.286242e-08, 
    -1.390616e-07, 2.670356e-08, -1.443948e-08, 2.27601e-10, -7.33155e-09, 
    2.299748e-08, 5.071001e-09, 1.530509e-08, 5.757704e-08, -1.894364e-09, 
    -1.61117e-08, 6.387756e-08, 1.469925e-08, 7.815231e-08, 2.545039e-08, 
    1.050512e-08, -3.237713e-08, -5.958839e-09, -1.102959e-07, 1.432796e-07, 
    9.681967e-08, -2.293825e-08, -1.84471e-07, -5.678016e-08, 2.292381e-09, 
    1.021317e-08, -6.234194e-08, -3.790191e-08, -3.186728e-08, -2.383878e-09, 
    1.249215e-08, -2.386663e-07, -5.828695e-08, 7.042151e-08, -3.25098e-08, 
    4.013145e-10, -1.364899e-07, -8.011385e-08, -4.32637e-07, 2.705335e-09, 
    6.595087e-09, 6.877769e-08, -1.949938e-07, 1.842836e-07, 8.243455e-08, 
    1.388377e-07, -7.446465e-08, -3.671312e-08, -2.983575e-08, -4.670937e-09, 
    8.760458e-08, 2.10722e-08, -1.614281e-07, -8.116103e-09, 1.635351e-08, 
    -3.01236e-09, -1.211463e-08, -5.419793e-09, -4.06616e-09, -4.678509e-08, 
    -2.89932e-07, -7.791864e-08, -1.81793e-07, -1.187332e-07, -5.201764e-08, 
    -4.44079e-08, -2.445984e-08, 6.921823e-09, -2.263484e-07, -3.448757e-07, 
    6.816663e-10, -6.02515e-08, 1.045308e-08, 1.691946e-07, -5.711627e-09, 
    3.537657e-07, -5.248513e-09, -3.580271e-08, -8.146355e-08, -1.688231e-08, 
    -1.599426e-08, -5.086351e-08, -7.215519e-09, -6.667385e-09, -4.39677e-08, 
    6.511698e-08, 1.442231e-08, -1.090848e-08, 1.264561e-08, -2.024774e-08, 
    -1.869262e-08, 5.598054e-09, 4.657022e-08, 9.440441e-09, -7.400558e-09, 
    2.428521e-09, -4.24042e-09, -6.104486e-10, 1.086214e-09, -2.675051e-08,
  1.013001e-08, 4.831446e-08, -3.670891e-09, -2.149903e-08, 1.552831e-08, 
    -8.61121e-10, 7.732353e-09, 1.147913e-08, -2.101154e-08, -5.622888e-08, 
    -8.537978e-08, -3.423719e-08, 7.248104e-10, -3.380791e-08, 2.457057e-09, 
    1.577023e-08, 9.56504e-08, 1.531498e-08, 1.644207e-07, 7.392202e-09, 
    -3.818906e-07, 1.969164e-08, -1.829898e-08, 7.930169e-09, 1.049131e-08, 
    4.17952e-08, 4.01688e-08, 1.940663e-08, 5.055284e-08, 4.494206e-08, 
    -1.404618e-08, 8.692751e-08, 7.811269e-08, 2.798776e-07, 4.214547e-08, 
    1.813163e-08, -9.803557e-10, -7.249199e-09, -1.050561e-07, 1.284915e-07, 
    6.31639e-08, -2.808605e-08, -1.917493e-07, -6.220912e-08, -3.148614e-09, 
    5.254094e-09, -2.712824e-08, -4.352063e-08, -2.253372e-08, -2.911776e-09, 
    1.149574e-08, -2.156435e-07, -4.2111e-08, 7.694624e-08, -3.560007e-08, 
    6.032792e-10, -1.098596e-07, 7.514128e-08, -4.915507e-07, 2.886509e-09, 
    6.468838e-09, 2.374748e-09, -1.1788e-07, 1.409201e-07, 1.081286e-07, 
    3.302415e-08, -8.17875e-08, -5.395935e-08, -6.638004e-09, -2.749914e-09, 
    7.806017e-08, 8.431073e-09, -8.122532e-08, -7.970868e-09, -2.078314e-08, 
    3.89781e-09, -1.880979e-08, -8.46245e-09, -5.577331e-09, -7.402087e-08, 
    -3.113204e-07, -4.65612e-08, -3.284044e-07, 1.325719e-08, -8.538456e-08, 
    2.668975e-08, -8.650375e-09, 1.894733e-08, -2.329185e-07, -3.625157e-07, 
    4.464084e-09, -6.36857e-08, 5.840832e-09, 1.363099e-07, -1.652398e-08, 
    4.215329e-07, -1.948871e-08, -2.079508e-08, -9.50883e-08, -1.419042e-08, 
    -2.506852e-09, -8.324172e-08, -1.156021e-08, -7.420226e-09, 
    -1.020365e-07, 6.48169e-08, -6.06604e-08, -1.874866e-09, -3.380518e-08, 
    -2.948781e-08, -3.576537e-08, 3.920491e-10, 3.955728e-08, 4.078044e-08, 
    -1.508562e-08, 1.747833e-09, -2.850314e-09, -6.541967e-11, 1.405517e-09, 
    -2.510211e-08,
  6.803418e-09, 6.375552e-08, 2.626217e-08, -2.232804e-08, 1.619338e-08, 
    1.291374e-08, 1.29167e-08, 1.304539e-08, -3.786738e-09, -1.909183e-08, 
    -5.731619e-08, -2.839403e-08, -1.121026e-08, -1.465139e-09, 2.031874e-08, 
    2.643243e-08, 9.18991e-08, 9.669867e-08, 6.152918e-08, -9.876857e-08, 
    -8.671833e-08, -9.982688e-08, -1.116263e-08, 9.955158e-09, -6.7418e-09, 
    6.238412e-08, 5.360238e-08, 2.151677e-08, 3.169845e-08, 8.340265e-08, 
    -7.6829e-09, 3.169185e-07, 7.91992e-08, 3.398855e-07, 3.949066e-08, 
    3.343195e-08, 1.802232e-08, -8.712036e-09, -1.045138e-07, 1.164877e-07, 
    4.126053e-08, -5.94253e-08, -1.707234e-07, -7.497098e-08, 4.604448e-08, 
    1.238374e-08, 6.458771e-08, -5.168332e-08, -1.442826e-08, -4.445837e-09, 
    1.04674e-08, -1.405224e-07, -1.017585e-08, 7.985201e-08, -3.660943e-08, 
    4.122285e-10, -7.669979e-08, 8.692666e-09, -7.484405e-07, -2.080147e-08, 
    -1.153751e-09, -1.300359e-07, -6.292186e-08, 8.8682e-08, 1.3823e-07, 
    -7.231785e-08, -7.402485e-08, -1.839737e-09, 6.266987e-10, -1.427054e-09, 
    5.849012e-08, 3.887692e-09, -3.868814e-08, -2.790017e-08, -5.207577e-08, 
    4.209198e-09, -7.816851e-09, -6.792533e-09, -5.626413e-09, -2.082818e-07, 
    -3.246697e-07, -7.814694e-09, -4.502483e-07, 1.962445e-08, -1.088184e-07, 
    -7.209763e-08, 3.5742e-07, 4.006478e-08, -2.187932e-07, -3.649536e-07, 
    -5.393474e-09, -6.220231e-08, 6.777867e-09, 1.291627e-07, -1.948473e-08, 
    5.069369e-07, -2.766318e-08, -2.960024e-08, -1.115242e-07, -1.102513e-08, 
    5.13154e-09, -8.348878e-08, -1.309242e-08, -1.533439e-08, -9.302238e-08, 
    5.040118e-08, -8.194201e-08, -3.429761e-09, -4.393809e-08, -4.577527e-08, 
    -4.370673e-08, -2.272924e-08, 1.620737e-08, 8.510477e-08, -1.037102e-08, 
    1.581225e-09, -8.496542e-09, -4.242651e-11, 1.687638e-09, -3.961901e-08,
  -8.504344e-10, 4.441728e-08, 1.119216e-07, 3.230809e-09, 7.437563e-09, 
    1.249504e-08, 1.418704e-08, 2.479908e-09, 9.464713e-09, 8.312725e-09, 
    -2.97843e-08, -1.07421e-08, -1.28436e-08, 5.201571e-09, 5.101111e-08, 
    4.95956e-08, 1.102191e-07, 9.35874e-08, -1.364695e-08, -1.597843e-07, 
    -1.038399e-08, -1.069934e-07, 3.603441e-07, 3.411281e-07, -5.432202e-08, 
    4.738416e-08, 4.084308e-08, 2.158123e-08, 2.381569e-09, 2.197834e-08, 
    3.097796e-09, 2.0832e-07, 5.714816e-08, 3.169825e-07, 1.137408e-08, 
    1.200895e-07, 2.474015e-08, -1.043476e-08, -1.272644e-07, 8.978738e-08, 
    7.931136e-08, -2.173758e-07, -1.381562e-07, -8.322215e-08, 2.258463e-08, 
    2.515657e-08, 4.094471e-08, -4.776183e-08, -1.246298e-08, -5.704059e-09, 
    9.35124e-09, -5.085673e-08, 1.709739e-08, 8.405819e-08, -3.793685e-08, 
    -2.096385e-10, -5.280168e-08, -5.976558e-08, -7.842002e-07, 
    -3.442696e-08, -2.753666e-09, -1.519128e-07, -3.41858e-08, 7.22374e-08, 
    1.701125e-07, 4.046689e-08, -6.039608e-08, -7.864344e-09, 4.073968e-10, 
    -4.456581e-09, 5.857015e-08, -2.202984e-08, 1.140819e-08, -7.002274e-08, 
    3.08966e-09, -3.057664e-09, 2.983555e-09, -8.394039e-09, -3.929104e-10, 
    -1.583788e-07, -3.063379e-07, -6.975375e-09, -5.177176e-07, 
    -1.295956e-08, -1.2753e-07, -1.627389e-07, 1.594285e-07, 3.299505e-08, 
    -2.005807e-07, -3.487171e-07, -3.801989e-08, -5.360076e-08, 7.110003e-09, 
    1.39208e-07, -2.429857e-08, 5.320325e-07, -5.516073e-08, 8.234196e-08, 
    -1.163499e-07, -2.538758e-08, -1.262725e-08, -4.382651e-08, 
    -1.308334e-08, -2.234263e-08, -3.652775e-08, 2.370081e-08, -7.25035e-08, 
    5.537117e-10, -3.652104e-08, -5.188741e-08, -2.751068e-08, -1.10558e-07, 
    8.678285e-10, 9.144452e-08, -4.211699e-09, 1.132366e-09, -1.661647e-09, 
    7.451462e-11, 1.874604e-09, -4.258766e-09,
  -2.854199e-08, 2.971092e-09, 1.414733e-07, 6.222399e-08, 2.48474e-09, 
    1.43018e-10, 1.062631e-08, -1.951867e-08, -1.130525e-08, 2.054844e-08, 
    -3.200739e-09, 2.448178e-08, 1.320996e-08, -9.920541e-09, 7.785866e-08, 
    6.368596e-08, 1.121798e-07, 3.448918e-08, -1.574588e-08, -2.261891e-08, 
    -2.825391e-08, -1.879903e-08, -3.378409e-08, 1.251533e-08, 5.102265e-10, 
    -6.350547e-09, 9.656105e-09, 2.390084e-08, -2.589627e-08, 8.908046e-09, 
    1.32884e-08, 7.953713e-08, -1.297622e-09, 3.412049e-07, -7.768449e-09, 
    4.339815e-07, 3.721566e-08, -1.029829e-08, -1.506935e-07, 3.466036e-08, 
    1.083584e-07, 2.311901e-07, -5.898522e-08, -8.154601e-08, -2.079605e-08, 
    2.52478e-08, 2.641349e-07, -3.766797e-08, -1.4856e-08, -7.589449e-09, 
    8.320285e-09, 2.679744e-07, 4.252258e-08, 8.690805e-08, -3.895202e-08, 
    -6.009486e-10, -3.95712e-08, 1.500487e-08, -5.374333e-07, -6.55416e-09, 
    -6.784148e-09, -7.837184e-08, -1.893886e-08, 3.982023e-08, 2.189485e-07, 
    3.717969e-08, -5.447214e-08, 1.38034e-08, -7.278231e-10, -1.723879e-08, 
    6.18079e-08, -3.052469e-08, 2.072375e-08, -7.369727e-08, 7.743599e-08, 
    2.323759e-09, 7.242932e-09, -3.839318e-09, 1.076484e-08, -9.116366e-08, 
    -2.768745e-07, -4.745397e-08, -5.468735e-07, -4.849107e-08, 
    -1.109247e-07, -9.423911e-08, -3.24103e-08, 2.14302e-08, -1.911193e-07, 
    -3.049046e-07, 4.957496e-08, -5.129077e-08, 3.234504e-09, 1.138429e-07, 
    -3.165928e-08, 2.512137e-07, -7.908634e-08, 3.722016e-08, -1.058752e-07, 
    -2.818665e-08, -4.945423e-08, -6.507645e-08, -1.129624e-08, 
    -2.540692e-08, 1.571152e-10, -1.325179e-08, -4.523395e-08, 7.423978e-09, 
    -3.583909e-08, -4.969274e-08, -1.507919e-08, -1.308269e-07, 
    -2.711931e-08, 3.132868e-08, -5.695051e-08, 4.329649e-10, 1.060528e-09, 
    1.447376e-10, 1.994266e-09, 1.395724e-07,
  -5.663316e-08, -3.745919e-08, 5.511976e-08, 4.639406e-08, -1.486347e-08, 
    -1.83033e-08, -2.099767e-08, -1.134898e-07, -6.397437e-08, 4.668431e-08, 
    -2.101916e-08, 2.165221e-07, -4.815871e-08, -2.856476e-07, 2.002167e-07, 
    7.515654e-08, 1.126222e-07, -1.31871e-09, 2.318713e-08, 1.635338e-07, 
    -7.157615e-08, -1.308155e-08, -4.848351e-08, -1.335678e-08, 3.276605e-07, 
    -5.180976e-08, -2.097823e-08, 2.352471e-08, -4.247346e-08, 9.559415e-09, 
    1.280983e-08, -4.723512e-08, -1.829477e-08, 4.594885e-07, -9.162989e-09, 
    3.125442e-07, 6.103953e-08, -8.324847e-09, -1.160203e-07, -2.956585e-09, 
    9.248905e-08, 1.295909e-07, -5.576788e-08, -7.286043e-08, -4.280986e-08, 
    2.077496e-08, 3.170057e-07, -9.695242e-09, -1.654952e-08, -8.529923e-09, 
    7.596427e-09, 5.186126e-08, 5.789908e-08, 8.536548e-08, -2.722342e-08, 
    -9.3587e-10, -3.847896e-08, 1.486729e-07, -2.976406e-07, 2.050672e-07, 
    1.208724e-08, -6.560259e-08, 5.014175e-08, 6.305561e-09, 2.383381e-07, 
    5.267054e-09, -3.270515e-08, 1.491514e-09, 2.546659e-08, -1.108248e-08, 
    6.318106e-08, 4.316519e-09, 4.414147e-08, -3.772124e-08, 9.934598e-08, 
    1.042366e-08, 1.207722e-08, -2.118577e-08, 1.95723e-08, -2.405574e-08, 
    -2.518862e-07, -5.83345e-08, -5.249054e-07, -6.230022e-08, -5.78404e-08, 
    1.579753e-08, -6.541819e-08, 1.535642e-08, -1.925882e-07, -2.552898e-07, 
    1.251927e-07, -4.457128e-08, 5.606353e-09, 6.790761e-08, -4.768953e-08, 
    1.661653e-07, -7.863981e-08, 3.515532e-08, -9.988599e-08, -1.656971e-08, 
    4.130868e-09, -7.539234e-08, -1.316101e-08, -1.946321e-08, 3.414453e-08, 
    -1.986933e-08, -1.127927e-08, 3.891103e-09, -3.861527e-08, -4.830764e-08, 
    -1.108646e-08, -5.460237e-08, -7.009083e-08, -5.475789e-08, 
    -4.425948e-08, -6.667847e-10, -7.591439e-10, -1.043645e-10, 2.208317e-09, 
    1.427563e-07,
  -8.991469e-08, -4.456956e-08, -3.055493e-08, -2.360935e-08, -3.249966e-08, 
    -3.585069e-08, -5.102561e-08, -1.480071e-07, -7.421522e-08, 1.195108e-07, 
    6.81614e-08, 2.161687e-08, -5.932611e-08, -1.614446e-07, 1.512649e-07, 
    8.254499e-08, 1.299127e-07, -6.676282e-08, 2.314357e-08, 1.387484e-07, 
    -1.358821e-07, 2.45094e-07, -1.91792e-08, -1.683254e-07, 1.168246e-07, 
    -9.305063e-08, 6.828486e-09, 1.771173e-08, -4.372578e-08, 4.647336e-08, 
    1.017634e-08, 4.124217e-08, -3.167179e-08, 2.868976e-07, 2.974048e-10, 
    2.193763e-07, 6.962973e-08, -6.554728e-09, -5.695188e-08, -9.693712e-09, 
    1.394169e-08, 7.337576e-09, -4.706243e-08, -6.223627e-08, -3.92572e-08, 
    5.290758e-09, 2.090179e-07, 2.091087e-08, -2.553156e-08, -8.064248e-09, 
    7.241198e-09, 1.025955e-08, 6.788514e-08, 8.143161e-08, -2.312091e-08, 
    -2.185629e-09, -3.519608e-08, 1.59212e-07, -5.901675e-07, -2.36447e-07, 
    1.793685e-07, 2.797492e-08, -1.038188e-09, 1.556259e-08, 2.311254e-07, 
    -1.85521e-08, -1.934222e-08, -2.753654e-08, -3.887862e-09, 1.7415e-08, 
    4.010735e-08, 5.381139e-08, 2.022762e-08, -3.697664e-08, 3.726114e-08, 
    1.073818e-08, 2.33108e-08, -3.007852e-08, 3.248411e-08, 1.498665e-08, 
    -2.379494e-07, -3.906629e-08, -4.474557e-07, -8.315465e-08, 1.661419e-08, 
    -1.667945e-08, -6.252276e-08, 1.043531e-08, -1.949451e-07, -2.297373e-07, 
    9.510609e-08, -4.012472e-08, 1.194968e-08, 2.932177e-08, -5.975448e-08, 
    1.010326e-07, -5.710645e-08, -4.816684e-08, -8.49252e-08, 3.4815e-09, 
    9.658993e-08, 5.195788e-08, -1.753125e-08, -1.209138e-08, 1.241754e-07, 
    -6.862592e-09, 9.026735e-11, -2.043043e-08, -4.36869e-08, -4.824142e-08, 
    -8.503321e-09, -1.547937e-08, -3.795458e-08, -2.018328e-08, 
    -7.124299e-09, -8.848019e-10, -2.989566e-09, -7.472636e-10, 2.492968e-09, 
    1.054377e-07,
  -2.161578e-07, -1.139392e-08, -5.316747e-08, -3.230616e-08, 1.508624e-08, 
    -4.874801e-08, -5.560742e-08, -2.048864e-09, -6.479968e-08, 3.022251e-09, 
    -4.430876e-08, -7.609492e-08, 1.566934e-07, 2.838578e-08, -3.971513e-08, 
    9.163573e-08, 1.825202e-07, -1.25006e-07, 4.268355e-08, 7.988024e-08, 
    -5.692186e-08, 1.119652e-07, 4.670665e-08, -7.225231e-08, -2.829797e-07, 
    1.856001e-07, -2.20507e-09, 1.666626e-08, -3.539117e-08, 1.184032e-07, 
    1.016724e-08, 7.229119e-09, -3.766218e-08, 1.185263e-07, 2.570323e-08, 
    2.996107e-07, 6.344862e-08, -5.23022e-09, -2.637921e-08, -2.535148e-08, 
    2.92031e-08, -3.093623e-08, -4.730038e-08, -5.165267e-08, -3.915898e-08, 
    -1.372223e-08, 8.31177e-08, 4.720562e-08, -3.454229e-08, -6.121454e-09, 
    7.115801e-09, -1.130695e-07, 6.197417e-08, 7.37809e-08, -2.569207e-08, 
    -9.320047e-10, -4.310323e-08, 2.769252e-08, -7.99147e-07, -1.147293e-07, 
    1.404169e-08, 2.937213e-08, -9.740165e-08, 2.669453e-08, 2.191997e-07, 
    1.640001e-08, -1.949275e-09, -2.988304e-08, -2.082606e-08, 1.618127e-08, 
    5.075663e-08, 1.0587e-07, -2.481329e-08, -1.021265e-07, -3.092193e-08, 
    1.60162e-09, 2.352016e-08, -2.352368e-08, 3.180028e-08, 8.8246e-09, 
    -2.238216e-07, -6.977031e-09, -3.554817e-07, -5.291736e-08, 3.142623e-08, 
    6.453752e-08, -6.196524e-08, 3.346941e-09, -1.797165e-07, -2.3655e-07, 
    -1.144247e-07, -2.854995e-08, 1.082287e-08, -8.634785e-09, -5.088191e-08, 
    4.789581e-08, -3.73298e-08, -6.623327e-08, -7.444419e-08, 1.750145e-08, 
    1.303638e-07, 1.404644e-07, -2.412077e-08, -8.618045e-09, 7.404697e-08, 
    2.523689e-08, -1.163198e-08, -4.334379e-08, -4.866365e-08, -5.10388e-08, 
    -8.282996e-09, -9.772975e-09, 3.553396e-09, 3.68118e-10, 1.38175e-09, 
    -3.433115e-10, -1.435836e-09, -1.016666e-09, 2.502617e-09, 5.351831e-08,
  -3.638232e-07, 2.286929e-07, 1.832135e-07, 9.089649e-08, 5.79422e-08, 
    -9.908399e-08, -5.580273e-08, -1.114566e-07, -8.030395e-08, 
    -1.338303e-07, -5.919492e-08, -7.285428e-08, -1.826246e-07, 1.396551e-07, 
    -1.896976e-07, 9.651497e-08, 1.942269e-07, -1.510567e-07, 6.868584e-08, 
    3.19834e-08, -6.726407e-08, -1.187534e-07, 7.162089e-08, -6.529672e-08, 
    -3.041328e-08, 3.430159e-08, 1.008754e-07, 1.441617e-08, -2.500565e-08, 
    9.769087e-08, 2.20366e-08, -5.515346e-08, -3.15456e-08, -1.247463e-08, 
    6.306277e-08, 2.595741e-07, 5.367095e-08, -4.433659e-09, 1.587421e-08, 
    -3.597914e-08, 1.215069e-08, 1.025285e-07, -2.814431e-08, -4.396065e-08, 
    -2.092202e-08, -2.290653e-08, 1.687232e-08, 6.422809e-08, -4.024221e-08, 
    -4.901658e-09, 7.251046e-09, -5.644699e-08, 5.068695e-08, 6.295383e-08, 
    -2.349003e-08, -7.747758e-11, -5.351626e-08, -6.400656e-08, 
    -7.048305e-07, -5.320443e-08, 2.754064e-09, -1.790454e-08, -1.03665e-07, 
    3.035757e-08, 1.960433e-07, 3.444609e-08, 1.520198e-08, -3.705065e-08, 
    2.89815e-08, 7.067342e-09, 5.255799e-08, 1.041872e-07, -4.225194e-08, 
    9.356427e-11, -3.889051e-08, -1.337469e-08, 2.993195e-08, -1.8571e-08, 
    1.126683e-08, -3.590515e-08, -2.145385e-07, 3.013756e-08, -2.883343e-07, 
    -4.576987e-08, -4.437197e-10, 1.776166e-07, -1.098283e-07, -1.33324e-08, 
    -1.778844e-07, -1.632737e-07, -8.073653e-08, -2.504478e-08, 6.284978e-09, 
    2.910039e-08, -3.871332e-08, 1.032708e-07, 1.788288e-08, -8.198026e-08, 
    -6.871369e-08, 2.325476e-08, 9.391908e-08, 1.696129e-07, -3.545009e-08, 
    -5.347566e-09, 6.469133e-08, -3.261835e-08, -4.213007e-09, -6.083928e-08, 
    -5.468507e-08, -5.501511e-08, -6.479581e-09, -7.880317e-09, 9.908717e-09, 
    6.879191e-10, 2.80113e-09, -3.125138e-10, -7.736247e-10, -2.281681e-09, 
    2.049106e-09, 9.489838e-08,
  -4.014036e-07, 7.178509e-07, 8.873722e-07, 2.887898e-07, 1.134367e-07, 
    -7.205233e-08, -7.486335e-08, -1.424734e-07, -6.005121e-08, 
    -7.687902e-08, -2.641548e-08, -5.089271e-08, -1.721173e-08, 2.523143e-08, 
    -1.618522e-07, 7.628768e-08, 1.649062e-07, -1.954191e-07, 4.400042e-08, 
    1.278933e-07, -1.207673e-07, -2.742274e-08, 4.541789e-08, 1.601347e-08, 
    -9.840846e-09, 7.722304e-08, 3.731088e-08, 1.380556e-08, -1.664444e-08, 
    1.0757e-07, 3.238756e-08, -1.084157e-07, -2.757736e-08, -1.125176e-07, 
    1.467737e-07, 2.955862e-07, 3.926703e-08, -3.411913e-09, 4.451067e-08, 
    -5.307275e-08, 8.819318e-08, -9.053338e-09, -6.981369e-08, -4.862622e-08, 
    -3.857167e-08, -1.846377e-08, -3.268474e-08, 7.130214e-08, -4.180876e-08, 
    -4.169337e-09, 7.596597e-09, -2.58799e-08, 3.765843e-08, 5.322711e-08, 
    -2.107626e-08, -1.184333e-09, -8.403015e-08, -1.397325e-07, -5.6589e-07, 
    -2.581959e-08, 1.288618e-08, -1.413446e-08, 2.153798e-07, 3.51959e-08, 
    1.897013e-07, 3.869559e-09, 2.592299e-08, -3.232708e-08, 5.962102e-08, 
    1.476815e-08, 1.592718e-08, 2.993033e-09, -6.319613e-08, 3.421951e-08, 
    8.475141e-09, -1.636306e-08, 2.940962e-08, -9.171259e-09, 2.348285e-09, 
    -8.757115e-08, -2.113595e-07, 1.371234e-08, -2.403166e-07, 1.249732e-07, 
    2.0176e-08, 1.143429e-07, -1.65956e-07, -6.035089e-08, -1.302658e-07, 
    -1.291502e-07, -4.555807e-08, -2.868696e-08, -5.337171e-09, 1.697078e-08, 
    -3.442722e-08, 2.124824e-07, 7.18964e-08, 2.622812e-08, -4.731919e-08, 
    2.091545e-08, 7.005724e-09, 6.872375e-08, -4.449388e-08, -6.006424e-09, 
    2.891466e-08, 1.244052e-08, -1.718945e-09, -7.465258e-08, -6.229368e-08, 
    -5.968661e-08, -5.360675e-09, -7.329845e-09, 1.144406e-08, 6.66887e-10, 
    3.744958e-09, -4.957879e-11, -1.018705e-09, -2.070003e-09, 1.37549e-09, 
    4.901142e-08,
  -7.321136e-07, 2.025167e-07, 5.885658e-07, 2.80243e-07, 1.017098e-07, 
    7.338485e-11, -4.445172e-08, -2.939652e-08, -6.714515e-09, 1.625693e-08, 
    1.932e-08, -6.714021e-08, 8.270092e-09, 6.922556e-08, -1.011989e-07, 
    4.470774e-08, 1.236862e-07, -1.37802e-07, 1.067529e-08, 1.853383e-07, 
    9.735061e-09, 4.678725e-09, 4.252792e-08, 3.040708e-08, -6.506468e-09, 
    2.835687e-07, 8.435961e-09, 1.131701e-08, -9.522694e-09, 1.503652e-07, 
    9.150824e-09, -2.260735e-07, -3.498923e-08, -1.222335e-07, 2.530215e-07, 
    6.751958e-08, 2.088931e-08, -2.058428e-09, 6.613874e-08, -5.757969e-08, 
    1.303231e-07, -1.905204e-08, -5.480058e-08, -4.965596e-08, -1.402776e-08, 
    1.230717e-09, -6.736781e-08, 8.824284e-08, -4.224299e-08, -1.854325e-09, 
    8.117254e-09, 9.254251e-08, 2.515193e-08, 4.149769e-08, -2.049764e-08, 
    -3.658442e-10, -1.239057e-07, -2.198483e-07, -4.31554e-07, -6.753585e-08, 
    1.113716e-08, 4.32222e-08, -4.571342e-08, 5.801681e-08, 1.740324e-07, 
    2.672499e-08, 2.703786e-08, -1.429777e-08, 7.750651e-08, 8.753602e-09, 
    -7.366026e-08, -1.280222e-08, -6.643239e-08, 5.959117e-08, -2.5416e-08, 
    -2.739893e-08, 4.431996e-09, -4.364372e-08, -3.708729e-09, -2.621454e-08, 
    -2.003789e-07, 2.282124e-09, -1.907036e-07, 2.293869e-07, 1.753637e-08, 
    7.932437e-08, -2.230649e-07, -1.279308e-07, 8.11653e-10, -1.077174e-07, 
    5.98863e-08, -3.44745e-08, -5.400963e-08, 4.038171e-08, -4.589396e-08, 
    2.723275e-07, 9.237006e-08, 1.591673e-09, -3.651525e-08, 1.49758e-08, 
    -2.54829e-10, 1.583935e-09, -2.201276e-08, -6.071232e-09, 1.180518e-08, 
    -8.484051e-09, -2.948411e-09, -8.665103e-08, -7.037835e-08, 
    -6.414649e-08, -4.903029e-09, -7.120377e-09, 1.291261e-08, 5.543939e-10, 
    3.588809e-09, 9.440213e-10, -1.34186e-09, -7.853771e-10, 1.015238e-09, 
    -1.059215e-08,
  -3.653223e-07, 4.104095e-11, -7.741789e-08, 8.812128e-08, 1.784491e-07, 
    1.786564e-07, 3.515754e-08, 6.927348e-08, 3.802609e-08, 1.900628e-08, 
    -7.245376e-09, 1.39537e-08, 9.508312e-09, 4.128856e-08, 4.22325e-08, 
    6.953599e-08, 8.321004e-08, -6.547458e-08, 2.213582e-09, 5.84381e-08, 
    5.31868e-08, 1.932256e-08, 4.076981e-08, 3.944876e-08, -7.403969e-09, 
    -2.611455e-08, 6.244022e-08, 1.216347e-08, -1.571448e-08, 4.059939e-08, 
    -5.520076e-08, -2.934636e-07, -4.202082e-08, 4.216145e-08, 2.31563e-08, 
    -2.140605e-07, 3.78983e-09, -1.134111e-09, 5.255754e-08, -5.237465e-08, 
    1.092035e-07, -2.257093e-08, -3.498911e-08, -3.281095e-08, -1.418061e-08, 
    -2.048512e-08, -9.645976e-08, 1.009561e-07, -2.155798e-08, 1.508745e-09, 
    8.799262e-09, 3.508848e-07, 1.232362e-08, 2.967406e-08, -2.011889e-08, 
    -2.13123e-09, -1.477073e-07, -2.798144e-07, -3.166717e-07, -2.846551e-08, 
    -9.886662e-09, 3.703383e-08, -4.440108e-08, 5.662337e-08, 1.385463e-07, 
    2.331899e-08, -3.894911e-10, 6.408277e-08, 9.301232e-08, 6.290406e-09, 
    -1.080723e-07, -1.094838e-08, -5.590664e-08, -3.695732e-09, 
    -3.303123e-08, -4.181948e-08, 1.068931e-07, -3.109537e-08, 2.344748e-09, 
    1.316494e-08, -1.890811e-07, 1.728615e-08, -1.44407e-07, 9.226596e-09, 
    -1.647288e-08, -1.203603e-08, -1.749366e-07, -9.164569e-08, 
    -6.338878e-08, -1.026978e-07, 6.185928e-09, -1.479223e-08, -1.772207e-08, 
    5.882441e-08, -7.925144e-08, 2.819091e-07, 9.483369e-08, 8.456232e-08, 
    -5.004824e-08, 5.7497e-08, 1.412025e-08, -4.583075e-08, -5.679862e-08, 
    -5.830898e-09, 1.312219e-08, -6.23553e-08, -9.921791e-09, -9.858525e-08, 
    -7.807432e-08, -6.861978e-08, -4.946514e-09, -6.94763e-09, 1.416845e-08, 
    4.183676e-10, 1.792387e-09, 1.275726e-09, -3.262144e-09, -2.828813e-10, 
    1.02078e-09, -1.799629e-08,
  -5.579074e-08, 2.081146e-08, -7.924308e-08, 1.259576e-08, 1.210418e-08, 
    -1.083833e-09, 3.098324e-08, 2.409882e-08, 4.16556e-08, 3.023962e-08, 
    4.33385e-08, 3.741189e-08, 1.730172e-08, 3.894689e-08, 6.717943e-08, 
    1.018977e-07, 4.496847e-08, 6.8215e-08, 5.368108e-09, 3.332622e-08, 
    2.674943e-08, 2.456858e-08, 3.876124e-08, 4.350596e-08, -1.026928e-08, 
    -2.470989e-08, 5.182841e-08, 3.857332e-08, -3.672045e-08, 1.391698e-07, 
    -4.829695e-08, -3.089804e-07, -3.243673e-08, -1.961951e-07, 1.154018e-08, 
    -2.705082e-07, -6.747404e-09, -9.757599e-10, -1.514879e-07, 
    -4.540018e-08, 4.905112e-08, -2.316739e-08, -3.867785e-08, -4.479135e-08, 
    -1.845984e-08, -3.162199e-10, -1.262123e-07, 1.103409e-07, 1.083848e-08, 
    3.708507e-09, 9.607433e-09, -4.706845e-08, 9.09131e-10, 2.098374e-08, 
    -1.988887e-08, -5.817867e-09, -1.229031e-07, -3.055729e-07, 
    -2.361958e-07, 6.431111e-08, -9.906273e-09, 3.72001e-08, -4.385589e-08, 
    5.101393e-08, 9.780875e-08, -5.701685e-08, -5.388637e-08, 1.03755e-07, 
    9.363504e-08, -5.096297e-09, -1.782577e-07, -8.755649e-09, -4.79094e-08, 
    -1.901469e-09, -3.579456e-08, 1.276192e-09, -2.813394e-08, -2.019218e-08, 
    -1.929754e-09, 2.972144e-07, -1.6366e-07, 1.1665e-08, -1.282169e-07, 
    9.234839e-09, -1.972847e-08, 3.45695e-08, -1.493028e-07, 2.358098e-08, 
    -6.488728e-08, -1.043578e-07, -8.464269e-09, -3.649291e-09, 2.958302e-09, 
    6.12726e-08, -1.715425e-07, 3.371194e-07, 8.112808e-08, -2.026758e-08, 
    -2.591418e-08, -8.167799e-09, -5.275695e-09, -6.185069e-08, -4.06587e-08, 
    -3.880629e-09, 1.410177e-08, -9.701176e-08, -1.785503e-08, -1.025133e-07, 
    -8.742853e-08, -7.324394e-08, -5.384493e-09, -6.903008e-09, 1.492657e-08, 
    2.818865e-10, 1.44945e-09, 1.692047e-09, -4.084299e-09, 1.065601e-10, 
    1.613344e-09, -1.892982e-08,
  -3.37468e-08, 2.986326e-08, -6.037499e-08, 7.070639e-09, -6.059736e-09, 
    2.992238e-10, 7.085873e-09, 2.294973e-08, 4.006029e-08, 3.871287e-08, 
    4.125036e-08, 3.797186e-08, 1.609374e-08, 3.381729e-08, 7.822746e-08, 
    1.156798e-07, 1.02114e-08, 2.066258e-09, 6.020571e-09, 2.755201e-08, 
    2.943966e-08, 2.633556e-08, 3.59139e-08, 4.607114e-08, -1.063268e-08, 
    -2.403954e-08, 1.648937e-08, 1.925468e-08, -8.360757e-09, -4.73683e-08, 
    8.022198e-09, -2.373533e-07, -1.603444e-07, -2.387205e-07, 8.360757e-09, 
    -2.804732e-07, -1.12716e-08, -1.347956e-09, -1.575911e-07, -4.130997e-08, 
    4.523277e-08, -2.415982e-08, -4.827029e-08, -5.135505e-08, 7.423478e-08, 
    1.17288e-07, -1.53158e-07, 1.169394e-07, 8.133519e-09, 5.250143e-09, 
    1.058785e-08, -1.006899e-07, -8.044048e-09, 1.501576e-08, -1.982251e-08, 
    -5.496304e-09, -8.534494e-08, -3.312823e-07, -1.828601e-07, 
    -7.184127e-09, -5.274842e-09, 3.609284e-08, -4.342405e-08, 6.925825e-08, 
    6.717519e-08, 5.311381e-08, -1.265792e-07, 4.743811e-08, 8.293819e-08, 
    -2.424781e-08, -1.502715e-07, -2.923116e-09, 5.084758e-09, -1.39471e-09, 
    -3.780606e-08, 6.462187e-09, -3.603705e-08, -8.573238e-09, -9.371393e-09, 
    2.492786e-07, -1.0751e-07, -1.894663e-08, -1.597954e-07, 8.467168e-09, 
    -1.994727e-08, 2.426509e-08, -1.251017e-07, 2.986712e-08, -7.232374e-08, 
    -1.085722e-07, -1.288095e-08, -2.422121e-09, 4.049696e-09, 6.458574e-08, 
    -1.03076e-07, 3.908425e-07, 6.250057e-08, 2.527668e-08, -2.202682e-08, 
    -1.935523e-08, -5.215497e-09, -6.696854e-08, -3.779743e-08, 
    -2.555964e-09, 6.364189e-09, -4.308981e-08, -2.088041e-08, -9.241035e-08, 
    -7.759991e-08, -7.538392e-08, -6.527216e-09, -6.851451e-09, 1.523222e-08, 
    3.485638e-10, 9.356427e-10, 1.296757e-09, -4.730481e-09, -4.082416e-09, 
    1.82321e-09, -1.707463e-08,
  -3.899981e-08, 3.275682e-08, -4.897538e-08, 5.211632e-09, -1.197486e-08, 
    -7.212293e-10, 3.912874e-08, 2.179581e-08, 3.928562e-08, 4.124604e-08, 
    4.099502e-08, 4.022445e-08, 1.42993e-08, 3.185164e-08, 8.565098e-08, 
    9.068859e-08, -7.414513e-11, -2.47278e-08, 6.866969e-09, 2.400225e-08, 
    2.857519e-08, 2.707361e-08, 3.186642e-08, 4.6384e-08, -1.20092e-08, 
    -2.464685e-08, 6.071105e-09, -9.86538e-08, -4.765411e-08, -5.2117e-08, 
    6.244591e-09, -2.130378e-07, -5.57468e-08, -2.722109e-07, 6.963546e-09, 
    -2.765942e-07, -1.3155e-08, -1.365294e-09, -7.082872e-08, -3.266835e-08, 
    3.692021e-08, -2.300249e-08, -3.0808e-08, -3.502046e-08, 1.075696e-07, 
    1.555975e-07, -1.737436e-07, 1.221279e-07, -2.315844e-09, 5.70337e-09, 
    1.174263e-08, -1.135284e-07, -1.381611e-08, 1.044295e-08, -1.9834e-08, 
    -5.714128e-09, -5.4471e-08, -3.48285e-07, -1.572829e-07, -9.385076e-09, 
    -6.959908e-09, 3.505966e-08, -4.311232e-08, 5.92619e-08, 6.770165e-08, 
    -3.985861e-09, -1.808535e-07, 7.742233e-08, -4.016397e-08, -2.765046e-08, 
    -9.350379e-08, -3.796458e-09, -1.760645e-08, -1.232138e-09, 
    -3.929221e-08, 7.556082e-09, -3.634219e-08, -1.430874e-08, -3.110856e-08, 
    2.138365e-07, -7.639312e-08, -3.671572e-08, -1.609978e-07, 7.822564e-09, 
    -1.972057e-08, -4.380718e-08, -9.969085e-08, 3.060427e-08, -8.057846e-08, 
    -1.105824e-07, -1.445551e-08, -1.999979e-09, 5.60135e-09, 4.841756e-08, 
    -7.741278e-08, 4.432792e-07, 6.814621e-08, 3.016453e-08, -3.350283e-08, 
    -2.167217e-08, -4.738467e-09, -6.836149e-08, -3.578903e-08, 
    -1.924889e-09, 1.235685e-08, -3.027617e-08, -1.209901e-08, -8.380493e-08, 
    -7.101335e-08, -6.699975e-08, -7.132257e-09, -6.607706e-09, 1.530611e-08, 
    3.221885e-10, -6.089977e-09, 2.811384e-09, -3.550241e-09, -1.359346e-08, 
    1.506393e-09, -1.313606e-08,
  -4.064992e-08, 3.339329e-08, -4.092789e-08, 3.583466e-09, -1.453651e-08, 
    -1.130473e-08, 3.757492e-08, 2.041787e-08, 3.850465e-08, 4.371321e-08, 
    4.066493e-08, 4.124303e-08, 1.459233e-08, 3.228575e-08, 8.880562e-08, 
    1.966872e-08, 1.484965e-09, -2.984535e-08, 7.658201e-09, 2.183521e-08, 
    2.776352e-08, 2.741598e-08, 2.883934e-08, 4.541408e-08, -1.586449e-08, 
    -2.271184e-08, 1.378788e-08, -1.055906e-08, -4.0609e-08, -3.823305e-08, 
    1.84599e-09, -2.581967e-07, -6.597571e-08, -2.651378e-07, 6.166204e-09, 
    -2.736569e-07, -1.351377e-08, -1.185612e-10, -2.279791e-08, 
    -2.741204e-08, 2.630878e-08, -2.048995e-08, -3.474156e-08, -1.892316e-08, 
    3.685039e-08, 1.426365e-07, -1.909667e-07, 1.256146e-07, -8.1974e-09, 
    4.977636e-09, 1.31693e-08, -1.195191e-07, -1.745502e-08, 6.88857e-09, 
    -1.980071e-08, -4.050946e-09, -4.241969e-08, -3.582181e-07, 
    -1.451744e-07, -9.573199e-09, -8.406857e-09, 3.663689e-08, -4.292536e-08, 
    5.518945e-08, 7.131449e-08, -1.070435e-08, -4.985583e-08, 9.00497e-08, 
    -5.126589e-08, -5.835489e-09, -4.94785e-08, -5.113463e-09, -3.449207e-08, 
    -5.749712e-10, -4.041188e-08, 1.030418e-08, -3.630588e-08, -1.780987e-08, 
    -2.704151e-08, 1.415665e-07, -4.488879e-08, -4.055995e-08, -1.584502e-07, 
    7.057622e-09, -1.94147e-08, -1.046247e-07, -7.770046e-08, 3.045005e-08, 
    -8.541558e-08, -1.110428e-07, -1.502946e-08, -7.069847e-10, 6.200139e-09, 
    3.872126e-08, -7.952673e-08, 4.857441e-07, 6.209835e-08, 3.296469e-08, 
    -3.36351e-08, -2.25035e-08, -4.394167e-09, -6.873076e-08, -3.526079e-08, 
    -3.486988e-10, 1.507971e-08, -2.611199e-08, 8.481663e-09, -8.267642e-08, 
    -6.976933e-08, -5.80572e-08, -5.524214e-09, -5.748404e-09, 1.421239e-08, 
    1.043077e-10, -2.659186e-08, 3.206878e-09, -4.744805e-09, -4.404299e-11, 
    2.747527e-10, -1.533834e-08,
  -4.142163e-08, 3.290887e-08, -3.56485e-08, 2.024706e-09, -1.579173e-08, 
    -1.464883e-08, 3.813699e-08, 2.011637e-08, 3.76204e-08, 4.607676e-08, 
    3.998395e-08, 4.171017e-08, 1.611983e-08, 3.311692e-08, 9.20632e-08, 
    -4.829052e-08, 2.274295e-09, -3.203832e-08, 8.728293e-09, 1.909865e-08, 
    2.632152e-08, 2.694975e-08, 2.658356e-08, 4.370571e-08, -1.949542e-08, 
    -2.568282e-08, -2.152603e-09, -1.975053e-08, -1.688392e-08, 
    -2.987741e-08, 8.405948e-09, -1.931722e-07, -8.958676e-08, -2.06572e-07, 
    5.424511e-09, -2.765723e-07, -1.332238e-08, -3.176126e-11, -5.309687e-09, 
    -2.537829e-08, 1.323679e-08, -1.76513e-08, -3.492937e-08, -1.503411e-08, 
    4.627793e-09, 1.075054e-07, -2.045527e-07, 1.272611e-07, -2.123598e-08, 
    6.096656e-09, 1.491939e-08, -1.225841e-07, -1.936879e-08, 4.606693e-09, 
    -1.98379e-08, -1.48475e-09, -3.606368e-08, -3.623825e-07, -1.396728e-07, 
    -9.397141e-09, -9.718917e-09, 3.797987e-08, -4.314353e-08, 5.266671e-08, 
    7.002151e-08, -5.302411e-09, 1.537745e-08, 9.960939e-08, -3.819304e-08, 
    1.536097e-08, -4.550594e-08, -8.479049e-09, -4.037878e-08, -9.328005e-11, 
    -4.151955e-08, 8.915151e-09, -3.604106e-08, -1.742856e-08, -3.120622e-08, 
    1.22665e-07, -2.474656e-08, -4.123709e-08, -1.539319e-07, 5.951449e-09, 
    -1.905761e-08, -1.142191e-07, -6.185502e-08, 2.990049e-08, -8.56882e-08, 
    -1.108291e-07, -1.455732e-08, 1.113211e-09, 6.345033e-09, 3.496798e-08, 
    -1.737163e-08, 5.12598e-07, 5.806404e-08, 3.386884e-08, -3.730617e-08, 
    -2.287799e-08, -3.830735e-09, -6.772419e-08, -3.397877e-08, 8.282086e-11, 
    1.697555e-08, -2.307257e-08, 5.298165e-08, -9.162244e-08, -7.238276e-08, 
    -5.1879e-08, -2.942613e-09, -3.29868e-09, 1.275174e-08, 2.94051e-10, 
    -5.242026e-08, -4.350704e-09, -4.866607e-09, 1.240963e-10, -3.278878e-09, 
    -1.90177e-08,
  -4.180123e-08, 3.157885e-08, -3.254883e-08, 4.834533e-10, -1.663142e-08, 
    -1.605571e-08, 4.175052e-08, 2.118753e-08, 3.667498e-08, 4.403825e-08, 
    4.119505e-08, 4.167731e-08, 1.482164e-08, 3.386248e-08, 9.304955e-08, 
    -4.43833e-08, 2.755371e-09, -3.370315e-08, 9.421541e-09, 1.642894e-08, 
    2.511302e-08, 2.660903e-08, 2.446706e-08, 4.20203e-08, -2.338805e-08, 
    -2.451731e-08, -1.004884e-08, -1.756638e-08, -6.543075e-09, -2.6799e-08, 
    -1.44974e-08, -1.917692e-07, -1.037748e-07, -1.67836e-07, 4.897117e-09, 
    -2.804558e-07, -1.289088e-08, -7.976695e-10, -2.483063e-08, 
    -2.195762e-08, 1.033959e-08, -1.578877e-08, -3.512721e-08, -7.231179e-09, 
    2.466436e-10, 8.830892e-08, -2.134998e-07, 1.269468e-07, -3.500128e-08, 
    4.569671e-09, 1.708928e-08, -1.237794e-07, -2.085733e-08, 4.616743e-09, 
    -1.986788e-08, -1.943363e-09, -2.867711e-08, -3.593208e-07, 
    -1.362802e-07, -9.048321e-09, -1.099914e-08, 3.825181e-08, -4.307725e-08, 
    5.142455e-08, 6.770962e-08, -3.580965e-09, 3.010626e-08, 1.012797e-07, 
    -4.422412e-08, 3.236988e-08, -4.138991e-08, -1.341681e-08, -3.39233e-08, 
    -4.371259e-11, -4.234512e-08, 7.42051e-09, -3.571303e-08, -1.629351e-08, 
    -2.969768e-08, 1.058332e-07, -1.460506e-08, -4.320088e-08, -1.515987e-07, 
    5.236132e-09, -1.855966e-08, -1.237451e-07, -4.483553e-08, 2.877488e-08, 
    -8.380921e-08, -1.058872e-07, -1.501331e-08, 3.056778e-09, 6.290719e-09, 
    2.749398e-08, 1.579753e-08, 5.348784e-07, 4.020288e-08, 3.418489e-08, 
    -3.750796e-08, -2.289647e-08, -3.061984e-09, -6.696209e-08, 
    -3.293611e-08, 1.051234e-09, 1.867426e-08, -2.041605e-08, 9.858815e-08, 
    -1.031776e-07, -7.511875e-08, -5.199075e-08, -2.847344e-09, 
    -1.001865e-09, 1.239181e-08, 4.93344e-10, -7.180955e-08, -4.867048e-10, 
    -6.109047e-09, 9.626145e-09, 1.319634e-09, -1.86796e-08,
  -4.177861e-08, 2.910411e-08, -3.191991e-08, -1.065985e-09, -1.736447e-08, 
    -1.66545e-08, 4.449652e-08, 2.300231e-08, 3.533768e-08, 4.195471e-08, 
    4.246277e-08, 4.087957e-08, 1.093639e-08, 3.404244e-08, 9.130321e-08, 
    4.374917e-08, 2.551133e-09, -3.404989e-08, 1.004278e-08, 1.366396e-08, 
    2.524035e-08, 2.621704e-08, 2.18626e-08, 4.028271e-08, -2.772634e-08, 
    -2.378505e-08, -1.308325e-08, -1.451843e-08, -7.382198e-09, 
    -2.106475e-08, -2.394307e-08, -1.900389e-07, -1.067094e-07, 
    -1.179013e-07, 4.528204e-09, -2.824126e-07, -1.305579e-08, -4.049099e-10, 
    -5.655141e-08, -2.061913e-08, 4.397776e-09, -1.380346e-08, -3.329234e-08, 
    -6.1129e-09, -9.36268e-10, 6.387671e-08, -2.13964e-07, 1.245468e-07, 
    -4.708671e-08, 6.504479e-09, 1.928149e-08, -1.233823e-07, -2.206752e-08, 
    4.748506e-09, -1.990003e-08, -6.741061e-10, -2.600422e-08, -3.49999e-07, 
    -1.402393e-07, -9.537672e-09, -1.241216e-08, 3.924112e-08, -4.237933e-08, 
    5.018068e-08, 6.637657e-08, -9.409291e-10, 3.391693e-08, 1.0501e-07, 
    -4.337159e-08, 4.564089e-08, -4.06306e-08, -1.102757e-08, -3.344593e-08, 
    5.974243e-11, -4.424221e-08, 7.51885e-09, -3.386369e-08, -1.549932e-08, 
    -2.965963e-08, 9.886122e-08, -1.202176e-08, -4.472616e-08, -1.500327e-07, 
    4.413721e-09, -1.76662e-08, -1.259817e-07, -3.412941e-08, 2.677388e-08, 
    -8.076772e-08, -9.89649e-08, -1.511734e-08, 3.022603e-09, 6.058201e-09, 
    9.530723e-10, 2.752546e-08, 5.421357e-07, 3.802035e-08, 3.247425e-08, 
    -3.668407e-08, -2.287819e-08, -1.972637e-09, -6.567711e-08, 
    -3.180978e-08, 1.221167e-09, 2.064377e-08, -1.708048e-08, 5.79966e-08, 
    -1.101319e-07, -7.665e-08, -5.405417e-08, -5.248523e-09, -1.412161e-09, 
    1.366487e-08, -3.701075e-10, -7.941145e-08, 4.009734e-11, -9.786575e-09, 
    4.565454e-09, 1.561784e-08, -1.554446e-08,
  -4.108341e-08, 2.326243e-08, -3.493966e-08, -3.216144e-09, -1.823202e-08, 
    -1.564257e-08, 4.5739e-08, 2.298492e-08, 3.24373e-08, 3.846009e-08, 
    4.099485e-08, 3.812198e-08, 7.929145e-09, 3.107124e-08, 8.551098e-08, 
    1.447493e-07, 1.361592e-09, -3.266433e-08, 1.072102e-08, 1.001268e-08, 
    2.558676e-08, 2.52914e-08, 1.718621e-08, 3.71727e-08, -3.161091e-08, 
    -2.349935e-08, -1.445795e-08, -1.14897e-08, -5.279048e-10, -2.265307e-08, 
    -2.351868e-08, -1.736742e-07, -1.118014e-07, -1.022964e-07, 4.338574e-09, 
    -2.790294e-07, -1.528758e-08, -1.627825e-09, -5.938006e-08, 
    -2.244874e-08, 3.865807e-09, -1.00402e-08, -4.052455e-08, -4.679919e-09, 
    -3.798903e-09, 3.649615e-08, -1.967021e-07, 1.196564e-07, -6.688621e-08, 
    7.279134e-09, 2.337455e-08, -1.198449e-07, -2.318555e-08, 1.434881e-08, 
    -1.988001e-08, 2.781917e-09, -2.886298e-08, -3.279912e-07, -1.300841e-07, 
    -9.942383e-09, -1.452014e-08, 4.201564e-08, -4.000566e-08, 4.681634e-08, 
    5.15677e-08, -1.753222e-09, 3.938618e-08, 9.469403e-08, -5.041176e-08, 
    4.848965e-08, -4.002419e-08, -1.410882e-08, -2.132828e-08, -1.290346e-11, 
    -4.349508e-08, 6.518519e-09, -3.241986e-08, -1.4184e-08, -3.429564e-08, 
    9.975935e-08, -9.418272e-09, -4.403392e-08, -1.4656e-07, 4.227275e-09, 
    -1.553002e-08, -1.229226e-07, -2.628127e-08, 2.226835e-08, -7.611189e-08, 
    -9.117497e-08, -1.130803e-08, 2.726562e-09, 5.452335e-09, -2.98474e-08, 
    3.032227e-08, 5.297351e-07, 3.339784e-08, 3.023405e-08, -3.443819e-08, 
    -2.176943e-08, 2.327738e-10, -6.256692e-08, -2.987485e-08, 5.990373e-10, 
    2.422161e-08, -1.049847e-08, 5.0251e-08, -1.133307e-07, -7.745376e-08, 
    -5.503927e-08, -6.34617e-09, -1.940805e-09, 8.88366e-09, 7.8673e-09, 
    -8.088301e-08, 1.411991e-10, -3.573334e-09, -1.106315e-11, 9.715791e-09, 
    -1.075711e-08,
  1.394873e-13, 4.817733e-13, 4.822437e-13, 1.093431e-13, -1.308238e-13, 
    -2.516544e-13, -4.172638e-13, -4.507576e-13, -5.374822e-14, 5.239709e-13, 
    5.173789e-13, -2.487903e-13, -1.75438e-13, 1.404567e-13, 2.087358e-13, 
    -4.38563e-14, 1.363051e-13, -8.859605e-13, -1.808729e-14, 2.937248e-13, 
    -6.339399e-13, -2.051598e-12, -6.176511e-13, 1.907519e-13, -1.972337e-13, 
    -2.023671e-13, -2.853297e-14, -4.666252e-14, -2.047144e-13, 
    -8.787892e-14, -3.282922e-14, -8.659212e-14, -1.810019e-13, 
    -2.203249e-13, -2.309398e-13, -1.567195e-13, 6.921187e-13, -8.376698e-12, 
    3.342206e-13, -4.28436e-14, -9.300015e-14, 1.961804e-13, -6.282116e-14, 
    2.096939e-13, 1.388971e-13, -6.720725e-14, 1.535511e-13, 1.760317e-13, 
    9.013826e-13, -1.703915e-12, -1.102639e-12, -8.474444e-13, 6.128156e-13, 
    2.667579e-13, 3.236966e-13, -1.030554e-12, 9.83086e-14, 1.133694e-13, 
    1.077264e-13, -2.415984e-12, 9.679154e-13, 5.623446e-13, 5.438354e-13, 
    -6.037319e-13, -1.33797e-12, -1.773415e-13, 9.786102e-14, 2.998368e-13, 
    1.26349e-13, 8.432185e-14, -4.590774e-14, 8.083427e-14, 9.496575e-14, 
    -1.689483e-13, 7.271642e-14, -5.532645e-13, 1.324049e-12, 1.102692e-13, 
    -3.343584e-12, -1.270301e-12, -7.38043e-13, -1.955431e-12, -7.214202e-13, 
    3.25143e-14, 3.334715e-15, 1.559346e-14, -1.285819e-13, 4.950993e-13, 
    -3.254672e-13, 8.347061e-13, -4.136404e-13, 7.403385e-13, -3.510679e-13, 
    -3.402521e-13, 1.258454e-13, 1.314354e-13, 2.807868e-13, -1.844883e-13, 
    -4.553758e-13, 8.67118e-13, -1.403543e-12, -6.275838e-14, -1.630987e-12, 
    2.570189e-12, 7.79627e-14, 3.329456e-13, 3.614518e-13, 9.235452e-13, 
    1.011472e-12, 5.386247e-13, 4.12226e-13, 3.421294e-14, 1.597464e-13, 
    1.609379e-13, 6.805529e-13, 5.28398e-13, -4.525896e-13, 2.543607e-13, 
    3.029892e-13, -1.650459e-12,
  -3.847336e-13, -3.579565e-13, -2.921442e-13, -2.956991e-13, -2.19165e-13, 
    -1.569005e-13, -1.231873e-13, -9.755259e-14, -2.477282e-13, 4.719848e-14, 
    -1.031352e-13, 1.623071e-14, -1.065375e-13, 4.096854e-13, 7.650694e-13, 
    1.123427e-13, 1.696539e-13, -1.806026e-13, -2.827716e-13, 7.139931e-14, 
    6.507278e-13, 1.495169e-12, 2.257614e-12, 1.784447e-14, 5.477993e-14, 
    1.974732e-13, 1.638812e-13, 1.842183e-13, 2.057181e-13, -6.543766e-14, 
    -1.368045e-13, -9.940712e-14, -1.27338e-14, -1.846652e-14, -8.525029e-14, 
    -7.377577e-14, -4.008012e-12, -1.473158e-13, -2.584142e-13, 3.255691e-13, 
    8.744482e-14, -2.432767e-13, -9.808285e-14, 1.694706e-13, 1.021432e-13, 
    7.75019e-13, -6.060218e-13, -5.082255e-13, 5.449175e-13, 1.128991e-12, 
    4.43131e-13, -4.958065e-13, 1.066786e-13, -6.63767e-12, 6.01495e-13, 
    -1.368338e-13, -1.022685e-13, -2.762304e-13, 1.308721e-12, 3.017109e-12, 
    3.668715e-13, -2.597644e-13, -3.244555e-14, 3.309422e-13, 5.306415e-14, 
    -6.545958e-13, -2.57894e-13, -1.355973e-13, 2.428062e-13, 4.067357e-13, 
    1.271963e-12, 2.202865e-14, 7.939977e-13, 4.362944e-13, -3.390576e-13, 
    -2.288139e-13, 4.50193e-13, -2.461348e-13, 3.589641e-12, -1.488971e-12, 
    1.04226e-13, -1.258624e-13, 7.555889e-13, 1.5702e-13, -5.232375e-13, 
    -4.777137e-13, 2.600907e-13, -6.086986e-13, -1.475996e-13, 1.055435e-12, 
    -3.683265e-13, -7.815839e-13, 8.578534e-13, 2.237095e-13, -2.516875e-13, 
    4.047602e-13, -2.54678e-13, 4.677173e-13, 7.581578e-13, 3.610757e-15, 
    -1.057435e-12, 3.985617e-13, -4.482389e-13, 3.535381e-13, -1.876537e-13, 
    -3.86138e-13, 1.234061e-13, -1.334019e-12, -4.680757e-13, -2.076049e-13, 
    -1.892624e-13, 9.172682e-14, 3.265054e-13, 4.599983e-13, 3.051041e-13, 
    -9.233469e-13, 3.823242e-15, 4.774026e-12, 2.096688e-13, -3.095792e-13,
  -1.305345e-13, -2.354505e-13, -1.516426e-13, -6.764034e-14, 5.080658e-14, 
    4.600487e-14, -7.510659e-14, -7.736867e-14, -2.326611e-13, -1.345313e-13, 
    -8.923418e-15, 9.450773e-14, -6.591949e-15, 1.733336e-13, 1.714046e-13, 
    2.382511e-13, 4.794318e-13, 7.673029e-14, 2.783017e-14, 4.797551e-14, 
    7.223111e-13, 7.563394e-13, 7.153583e-13, -2.496614e-14, 1.084827e-13, 
    -1.067063e-13, -3.552159e-13, -1.007805e-13, -1.38195e-13, -1.030703e-13, 
    -1.647432e-13, -2.22794e-13, 1.139089e-13, 6.379619e-14, -4.157785e-14, 
    -3.724798e-14, -1.54599e-12, -1.176443e-12, -1.142142e-13, 1.790151e-13, 
    -3.943235e-13, 6.429579e-14, -2.148455e-13, 2.312245e-13, 2.280259e-13, 
    5.088152e-13, -1.680753e-12, -8.371359e-13, -1.363482e-12, -2.912115e-13, 
    -1.110223e-16, -1.683653e-13, -6.458972e-13, -5.415188e-12, 1.669838e-13, 
    1.721713e-12, 1.459111e-13, -1.036439e-12, 5.899045e-13, -9.922965e-14, 
    2.863543e-13, 1.270789e-13, -7.049916e-14, 5.75473e-13, 1.565942e-13, 
    5.613565e-14, -1.617456e-13, -2.614575e-14, -1.657285e-13, -2.338685e-13, 
    1.933079e-12, 1.905281e-13, -7.130407e-13, 9.23317e-13, 3.664874e-13, 
    -2.956246e-13, -1.464124e-13, 1.128635e-12, 2.145553e-12, 2.608885e-13, 
    3.436973e-13, -4.529571e-14, -3.061926e-13, 6.350614e-13, 9.079959e-13, 
    -4.38094e-13, 9.567347e-14, 7.601836e-13, 3.089783e-13, -4.437839e-13, 
    -1.741662e-14, -3.594236e-13, 2.139608e-13, -1.002061e-12, 1.164069e-13, 
    -1.389236e-13, -7.42037e-13, 7.810419e-14, 5.349748e-13, 4.336032e-13, 
    -6.280948e-13, 2.607029e-14, 1.69335e-14, -6.791442e-14, -1.025e-12, 
    2.830097e-13, 3.75644e-13, 7.837619e-13, 8.388151e-13, 7.141648e-13, 
    1.050021e-12, 2.639833e-13, 1.85893e-13, -9.552081e-14, 8.337775e-13, 
    2.475076e-13, 1.860862e-11, 2.586256e-14, -1.024277e-12, -1.089989e-12,
  -1.603578e-13, -2.122469e-13, -1.959266e-13, -1.622313e-13, -1.362938e-13, 
    -8.12822e-14, -4.61714e-14, -8.869294e-14, 1.101202e-13, 4.505146e-13, 
    6.767087e-13, -1.807859e-13, -1.49547e-13, 1.018075e-13, 3.382711e-13, 
    6.027678e-14, 5.546119e-14, 3.300832e-14, 3.366231e-14, -3.891193e-13, 
    1.183637e-13, 5.623974e-13, 4.672512e-13, -2.300521e-13, -2.053635e-13, 
    -4.309608e-13, -3.354816e-13, 4.834466e-13, 8.477941e-14, 2.766953e-13, 
    3.469447e-13, 2.525341e-13, 4.425627e-13, 4.175826e-14, -8.733292e-14, 
    -5.187517e-14, -1.013356e-13, -1.56518e-12, -1.90542e-13, 3.23741e-14, 
    5.714318e-14, -3.455847e-13, -6.442277e-13, 2.847288e-14, 2.151196e-13, 
    1.351461e-12, 2.921968e-14, -1.519097e-12, 6.080692e-14, 1.465191e-11, 
    1.222258e-12, -7.418649e-13, -1.683599e-12, 2.202544e-13, -1.093039e-13, 
    1.647724e-12, 2.451817e-12, -1.418748e-12, 5.214884e-13, -1.25277e-12, 
    5.50851e-13, -1.943307e-13, 6.48398e-13, 2.654543e-14, -1.422362e-13, 
    -8.867074e-13, -6.361994e-13, -1.139436e-12, -6.887962e-13, -3.44974e-13, 
    2.026476e-12, 1.048606e-13, 2.170625e-13, -6.938894e-17, -4.444015e-13, 
    -1.702735e-12, -6.296508e-13, 3.299576e-12, -2.060365e-11, 5.277723e-14, 
    5.513923e-13, 1.043191e-12, 1.209449e-13, -2.017553e-13, -1.479372e-14, 
    2.125244e-13, -7.790296e-13, -3.107237e-13, -1.04972e-12, -7.297843e-13, 
    9.994783e-14, -9.640649e-13, 9.763163e-13, 2.982015e-12, 1.923461e-14, 
    -2.419814e-13, 2.9029e-13, -2.168543e-13, -1.082551e-12, -6.692591e-13, 
    -8.418544e-13, -3.011064e-13, 5.830267e-13, -1.080218e-12, -1.911249e-13, 
    4.336392e-13, 7.687184e-13, 8.318485e-13, 9.298118e-13, 9.411083e-13, 
    8.392176e-13, 5.247053e-13, 2.273043e-13, -4.460321e-14, 5.341561e-14, 
    2.224901e-12, 6.860417e-12, -9.995998e-12, 2.179324e-13, 3.56451e-13,
  -4.989065e-14, -1.75096e-13, -1.978279e-13, -2.079864e-13, -1.464801e-13, 
    -1.901118e-13, -3.242545e-13, -3.91423e-13, -5.230677e-13, 9.762885e-13, 
    8.597428e-13, -1.044997e-14, -5.43135e-13, -4.51722e-14, 8.167078e-14, 
    2.399192e-14, -4.056477e-14, -2.730455e-13, -1.941398e-13, -6.702278e-13, 
    -1.086894e-12, -4.401063e-13, 8.139184e-13, -9.174606e-14, -7.931156e-14, 
    -3.593653e-13, -2.985112e-14, -1.150052e-13, -2.31079e-13, -6.371709e-13, 
    -1.025777e-12, 7.939899e-13, 6.149664e-13, 4.876516e-13, -1.181708e-12, 
    -1.578321e-13, 3.314016e-14, 3.294927e-12, 6.163819e-13, -1.451503e-12, 
    1.207914e-12, -1.186412e-13, -4.957701e-13, -2.719283e-13, 4.277537e-12, 
    6.838557e-13, 1.726674e-13, 2.947365e-12, 1.986164e-12, 2.113864e-11, 
    1.849767e-12, -3.236703e-12, 1.546718e-12, -7.223028e-13, 9.098209e-14, 
    1.882244e-13, -9.394291e-13, 2.923078e-13, 6.018242e-14, -1.094666e-12, 
    -2.80484e-13, -4.350825e-13, -6.903228e-13, -1.040362e-13, -2.978146e-13, 
    2.273876e-13, -5.494216e-14, 1.160322e-13, 7.919637e-13, 2.669906e-12, 
    3.84956e-13, -2.072925e-13, 5.99007e-13, 7.779472e-13, -5.431155e-13, 
    -1.502395e-12, 1.935768e-12, -1.330068e-12, 2.712225e-12, 4.252848e-13, 
    1.196473e-12, 1.000373e-12, 1.191686e-13, -1.053616e-12, -1.999095e-13, 
    1.869754e-13, -1.913608e-13, -1.022474e-12, 5.69998e-13, -2.324779e-12, 
    -4.815731e-13, 4.493489e-13, 3.383752e-13, 1.182884e-12, 2.635253e-13, 
    8.288559e-12, 4.985748e-12, -4.279771e-13, -5.158998e-12, 6.835282e-13, 
    -1.902936e-12, 5.665433e-14, 9.579143e-13, -1.845338e-12, -4.713313e-13, 
    1.030703e-13, 1.421224e-13, 2.316064e-13, 5.212358e-13, 3.038264e-13, 
    1.796202e-13, 3.231165e-13, -3.298889e-13, -1.031536e-13, -9.820894e-13, 
    1.531098e-12, 9.508908e-12, -1.425825e-11, -4.803016e-13, -7.367718e-14,
  -1.513234e-13, -4.357625e-13, -5.814793e-13, -6.195322e-13, -7.665812e-13, 
    -7.119305e-13, -3.174683e-13, 6.503686e-13, 6.264433e-13, 2.569611e-13, 
    -4.650724e-13, -7.203405e-13, 9.527656e-13, 2.44077e-12, 2.804701e-13, 
    2.571582e-13, -8.394396e-13, -6.911277e-13, -1.700029e-15, -6.374345e-13, 
    -1.538353e-12, -1.700029e-13, 7.941148e-13, 6.292189e-13, -1.397771e-13, 
    8.230361e-13, -2.749467e-13, -3.615719e-13, 3.306244e-13, -6.798728e-13, 
    -1.86734e-12, 3.218814e-13, -1.525391e-12, -7.408518e-13, -1.622674e-12, 
    3.795575e-13, -3.566869e-14, 3.367383e-12, 1.087075e-12, -1.215694e-14, 
    -1.084799e-13, -9.904161e-12, -7.052067e-13, -1.113727e-13, 3.679307e-12, 
    2.873035e-12, 4.217043e-13, -4.028791e-13, 3.220752e-12, 1.012669e-11, 
    6.178252e-13, -1.487088e-12, -3.869405e-14, 5.614009e-12, 6.930859e-13, 
    9.109657e-13, 2.009309e-12, 2.909783e-13, 2.60971e-12, 2.775086e-12, 
    1.396189e-12, -3.060469e-12, -1.349365e-12, -2.130962e-13, -7.479573e-13, 
    5.304923e-13, -5.598022e-13, -2.555095e-12, -3.857803e-12, 4.033773e-12, 
    -1.091544e-12, -1.057765e-12, 1.249001e-12, -1.029538e-12, 3.051615e-13, 
    -1.833311e-12, 3.079828e-14, -4.614642e-13, -5.202221e-12, -3.760381e-12, 
    1.028025e-12, -1.515653e-12, -1.41484e-13, 5.648537e-13, 1.916522e-13, 
    5.046075e-12, 3.174683e-13, -7.691348e-13, -2.754692e-12, 3.422554e-12, 
    -9.791057e-13, -3.412104e-13, -8.541085e-13, 2.477907e-13, 3.755329e-14, 
    2.338013e-12, -8.574641e-13, -9.728329e-14, 3.636813e-13, -1.824152e-13, 
    -6.214751e-13, 2.208882e-12, 5.235812e-13, -6.072727e-12, -4.472811e-13, 
    -1.183498e-13, -2.084444e-14, 2.885747e-13, 5.663248e-13, 2.708112e-13, 
    -4.727607e-13, 5.180578e-13, -2.051692e-13, 1.080802e-13, 1.261935e-12, 
    1.335482e-12, 5.273386e-13, 1.083267e-12, 5.461395e-13, -2.205153e-12,
  -7.562839e-13, 2.125522e-13, 2.163825e-13, 4.526934e-13, 2.305656e-12, 
    5.995759e-12, 4.417022e-12, 1.088019e-12, 2.569833e-12, 3.669842e-12, 
    3.344269e-12, -2.764455e-14, 5.117573e-13, 3.846423e-12, 1.367134e-11, 
    1.802725e-13, -2.15199e-12, 1.273981e-12, -1.796112e-12, -1.662614e-12, 
    -5.538348e-13, 8.931744e-14, -5.815903e-13, -9.094392e-13, 3.292366e-13, 
    4.172385e-12, 9.114931e-13, 1.17556e-12, -2.751688e-12, -4.857781e-12, 
    6.573631e-13, 4.032885e-12, 2.08461e-12, -2.302603e-12, -4.934497e-12, 
    -4.071743e-12, 6.064149e-13, -4.932096e-13, -1.806888e-13, 2.661649e-12, 
    4.360401e-13, -3.210432e-12, -2.010753e-12, 6.507104e-13, 6.126544e-12, 
    4.908796e-12, 2.127326e-12, -5.600659e-13, 5.953893e-12, 5.338469e-12, 
    3.28032e-12, -3.003153e-14, -1.686151e-13, 8.568401e-12, 1.171342e-12, 
    1.078027e-12, 1.197709e-12, 1.277661e-12, 4.485429e-12, 4.871874e-12, 
    5.545453e-12, -3.468725e-12, -4.121592e-12, -8.60223e-13, -1.418143e-12, 
    -4.023115e-12, -1.158224e-11, 6.297352e-12, 7.594425e-12, 2.031675e-11, 
    -3.669287e-12, 5.0977e-12, -1.335487e-12, -4.891088e-13, -4.64212e-13, 
    -1.365241e-12, -1.016617e-13, 8.96061e-13, -7.48214e-12, -4.933998e-12, 
    2.508771e-12, 4.263527e-12, -3.756717e-13, 3.112566e-12, -7.190915e-13, 
    7.045531e-12, 5.770218e-12, -2.504663e-13, 8.651517e-13, 3.179679e-13, 
    1.082967e-12, -1.095579e-12, -6.564194e-14, -3.765022e-12, 3.825162e-12, 
    -8.740614e-12, -2.332579e-13, 5.181411e-13, 5.242973e-12, 1.079126e-12, 
    1.775302e-12, 2.800205e-12, -1.020753e-12, -5.020201e-11, -7.84206e-13, 
    1.881828e-13, -9.212076e-13, -2.463585e-13, -5.720979e-13, -1.004641e-12, 
    -1.696976e-12, -4.624634e-13, -9.174883e-13, 2.747247e-13, -2.910006e-12, 
    8.493595e-13, 1.566525e-13, 4.993991e-13, 3.610584e-13, -2.797651e-12,
  -6.555867e-14, 1.21092e-12, 1.21908e-12, 3.712031e-12, 6.221357e-12, 
    1.863953e-12, 2.993938e-12, -1.058265e-12, -3.924028e-12, -3.757994e-12, 
    -6.305956e-12, 6.227241e-12, 1.540823e-12, 5.433209e-12, 5.394574e-13, 
    1.725681e-12, 2.942729e-12, -5.3407e-12, -3.862119e-12, 3.183231e-12, 
    2.306544e-12, 8.770762e-15, -2.393086e-13, -4.286016e-13, 7.222667e-12, 
    9.560186e-12, -2.41418e-12, -4.039991e-12, -1.387612e-12, -8.507195e-12, 
    1.301792e-12, 5.341394e-12, 9.820644e-12, -2.584877e-12, -3.662959e-12, 
    -1.391109e-13, -5.145606e-13, 8.420209e-13, 5.07594e-13, -1.038031e-12, 
    -7.137358e-12, 3.641754e-12, 2.688905e-12, 6.829069e-13, 4.400424e-12, 
    3.542944e-12, 4.027056e-12, -2.471356e-13, 2.083589e-12, 7.522802e-13, 
    5.757422e-12, 1.612099e-12, 3.78586e-15, 2.36422e-13, 5.716261e-13, 
    5.250245e-13, 1.36724e-12, 4.056161e-12, -1.461448e-12, 4.216801e-12, 
    3.053335e-12, 5.499545e-12, -2.808087e-12, 6.25553e-12, 3.200684e-12, 
    -8.019085e-12, -2.560829e-11, 1.061984e-12, 2.923917e-11, -1.876499e-12, 
    -4.949929e-13, -4.931e-12, -5.069278e-12, -5.646039e-13, -3.371758e-12, 
    -6.462053e-13, -1.844774e-13, 6.90184e-13, -3.124112e-12, 1.422029e-12, 
    5.063394e-12, 5.081265e-12, 2.650186e-12, -2.307043e-13, -2.416956e-13, 
    1.272316e-12, 1.773692e-12, 1.387945e-12, 2.126385e-12, -4.088119e-13, 
    3.194112e-13, 8.539836e-13, 4.816009e-13, 8.329671e-13, 1.847411e-12, 
    -1.295188e-11, -4.499046e-12, -1.003575e-11, 5.258849e-12, 2.15733e-12, 
    -4.372946e-12, 2.914835e-12, -5.570024e-13, -5.474743e-11, -7.484569e-13, 
    -3.43725e-13, -1.447509e-12, -7.110423e-13, -1.975253e-12, -1.732225e-12, 
    -2.355283e-12, -4.835521e-12, -7.815359e-12, -4.446776e-12, 
    -1.651457e-13, 7.743806e-14, -2.159661e-13, -1.267139e-12, -5.384235e-14, 
    5.977718e-12,
  3.642683e-12, 1.73693e-12, 4.275344e-12, 3.545428e-12, -5.344072e-12, 
    -5.720993e-12, -1.302715e-11, -1.566483e-12, 7.956651e-11, 3.524191e-11, 
    9.372364e-13, 2.708431e-12, 6.370876e-13, -2.746262e-12, -4.248171e-12, 
    4.854742e-12, 1.463804e-12, -1.24548e-11, 5.864684e-13, 2.637376e-12, 
    1.191686e-13, -3.844106e-12, -8.577541e-12, -1.238894e-11, 2.842934e-12, 
    -1.917584e-11, -1.847041e-11, -1.891444e-11, -2.194751e-11, 
    -1.633485e-12, -5.160455e-13, -9.465387e-12, -1.894943e-12, 
    -5.590112e-13, 2.201699e-11, -2.931462e-11, -6.11429e-12, 1.694818e-12, 
    4.433341e-11, 1.275416e-12, 1.3513e-11, 1.207187e-12, 9.848511e-13, 
    -2.73592e-12, 3.021347e-12, 3.82587e-12, 5.881115e-12, -7.450984e-13, 
    5.128317e-12, 2.441367e-12, 3.450878e-12, -4.170692e-13, -3.548356e-13, 
    3.491624e-13, 3.911316e-13, 6.404738e-13, -1.865522e-12, 6.76191e-12, 
    -8.394868e-13, 2.321402e-11, -7.894477e-12, 4.623843e-12, -5.650619e-13, 
    2.302444e-12, -1.18682e-12, -1.046134e-10, 5.434583e-12, -1.644365e-12, 
    8.912968e-12, 1.264364e-12, -3.07844e-12, 2.560036e-13, 1.047926e-12, 
    -1.312252e-11, -6.340381e-12, -2.409808e-12, -3.41005e-13, -7.345513e-14, 
    6.500797e-12, 1.013564e-12, 1.049412e-11, -5.21177e-11, 3.135339e-12, 
    -5.203962e-12, -5.354175e-12, -2.750369e-12, -1.826941e-12, 
    -1.085006e-11, -1.108801e-12, 1.081621e-12, 1.121145e-12, -5.830217e-12, 
    -1.651596e-13, 2.234088e-12, -2.556025e-12, -8.656778e-12, -1.184954e-11, 
    1.777416e-11, -1.163972e-12, 2.285846e-12, -8.898618e-12, 2.229755e-12, 
    2.483812e-13, -2.767437e-11, 2.746234e-12, 8.803375e-13, -2.154235e-12, 
    -5.325976e-12, -7.826198e-12, 7.682605e-13, -5.713444e-12, -1.011809e-11, 
    -1.163182e-11, -6.67634e-12, 7.355713e-12, 1.349504e-13, -7.910339e-15, 
    -2.097001e-12, 4.277828e-14, 5.413212e-12,
  -7.204015e-12, -2.849387e-12, -7.673306e-13, 4.135192e-12, 6.51762e-12, 
    -3.085421e-12, 3.496176e-11, 1.236595e-10, -1.446533e-10, -1.43348e-10, 
    4.732381e-12, -6.902201e-12, -1.526501e-11, 1.204692e-11, 1.832423e-13, 
    1.924105e-12, -1.128764e-12, -9.453632e-12, -2.530455e-12, 1.900646e-12, 
    -6.331491e-12, 4.267087e-12, 1.70805e-11, -3.062334e-11, 1.557199e-12, 
    1.281936e-11, -1.88039e-11, -9.447554e-12, 3.756273e-12, -4.207779e-11, 
    2.523631e-11, -9.754308e-12, -1.516676e-12, -7.278456e-12, 5.036443e-11, 
    -4.725109e-13, -1.121184e-11, 1.417907e-12, 1.189548e-12, 5.366674e-12, 
    7.826372e-12, -1.451839e-12, 1.426984e-12, -2.961568e-12, 1.829092e-12, 
    6.301404e-12, 6.167428e-12, -5.607598e-13, 7.385115e-12, 3.919878e-12, 
    9.150944e-13, -3.522738e-12, -1.054634e-12, 1.382761e-12, 1.06147e-13, 
    8.010814e-13, -2.349848e-11, 8.689766e-12, -1.645423e-12, 2.641769e-11, 
    -2.430972e-11, 9.215795e-12, 1.068978e-11, -8.903211e-13, -6.222622e-12, 
    -5.759282e-11, -1.067424e-12, 2.931494e-11, 3.788858e-12, 1.756884e-11, 
    -1.577721e-11, -3.061051e-12, 9.522938e-12, -8.685386e-12, -7.938538e-13, 
    -6.57685e-12, -5.588932e-13, 1.647474e-12, 7.035263e-12, 9.652168e-12, 
    6.41534e-12, -7.228992e-11, 1.76692e-13, 3.3683e-11, -1.565931e-11, 
    -9.069245e-12, -4.280354e-12, -1.084982e-11, -3.744704e-12, 2.457839e-12, 
    -9.904855e-13, -1.370477e-11, -7.693984e-13, 7.444044e-15, -1.522948e-12, 
    2.68785e-13, -6.379552e-12, -3.949546e-11, -1.04422e-12, 5.619949e-14, 
    -8.132717e-12, -2.130195e-11, -1.330221e-13, 6.692098e-12, 5.287104e-12, 
    5.796474e-12, 6.221301e-12, -3.343492e-12, -9.800716e-12, 4.57373e-12, 
    -1.337103e-11, -1.385597e-11, 3.705369e-13, 3.906209e-12, 6.039502e-12, 
    1.539879e-14, 8.856804e-14, -2.598432e-12, 3.03594e-13, 1.056299e-11,
  -3.409339e-11, 4.831135e-12, 6.786016e-12, 1.816092e-11, 2.912315e-11, 
    7.596213e-11, 1.174973e-10, 2.911427e-11, -5.578538e-11, 1.198586e-11, 
    -1.008649e-11, -6.118661e-12, -1.17617e-11, -5.687784e-12, -9.070744e-12, 
    1.688716e-12, -2.871681e-12, -4.079737e-12, -3.384196e-12, 4.978129e-12, 
    3.34599e-12, 1.72119e-11, 3.661405e-11, -7.908563e-12, 4.217837e-11, 
    -3.206069e-11, -1.946121e-11, -2.083334e-12, 1.677436e-12, -1.416778e-11, 
    1.358358e-11, -4.469503e-11, 3.739475e-11, -1.020439e-11, -1.903389e-11, 
    -3.193013e-11, -2.874567e-12, 8.088669e-13, -1.224809e-11, 6.685863e-12, 
    -6.929857e-12, 9.137469e-12, 3.977735e-12, -1.576746e-12, 3.460565e-12, 
    -1.102862e-11, 5.000333e-12, 2.025519e-12, 4.984946e-12, 7.019524e-13, 
    5.981465e-13, -2.017708e-11, -8.162027e-13, 8.310019e-13, 3.581024e-14, 
    2.279843e-13, 1.819489e-11, 7.681955e-12, -3.782141e-12, 6.250001e-11, 
    -2.518608e-11, -1.034728e-13, -1.994072e-12, -3.640532e-12, 
    -5.873879e-12, -1.421711e-10, -1.197009e-11, 9.189138e-11, 2.157008e-11, 
    3.080536e-12, -3.672507e-11, -2.150047e-11, 4.624079e-12, 6.080803e-12, 
    5.606382e-12, -5.293987e-12, -6.583345e-13, 6.280393e-12, -1.006584e-13, 
    8.425372e-12, 3.04895e-12, -1.326103e-11, -4.407585e-14, 4.661838e-11, 
    8.832046e-12, 1.094791e-11, -1.360275e-10, -8.126944e-12, -2.036768e-12, 
    1.787737e-12, 9.200529e-12, -1.327391e-11, -1.484951e-12, 1.046174e-12, 
    -4.70014e-11, -8.039347e-13, -3.745271e-12, 4.536271e-11, -6.587952e-12, 
    -3.293121e-12, -1.788691e-11, -3.677395e-11, 4.570858e-13, 1.151349e-11, 
    -4.198975e-12, -1.723721e-11, -1.263833e-11, 1.303413e-11, 4.336864e-12, 
    8.48932e-12, -8.411161e-12, -6.955214e-12, -9.365841e-13, 3.99536e-12, 
    3.420264e-12, 3.819167e-15, 3.185924e-13, -1.671892e-12, 1.009372e-11, 
    6.584955e-12,
  -1.786349e-12, -1.836553e-11, 2.104916e-11, 6.781131e-11, 1.519183e-10, 
    1.671558e-10, 5.946954e-11, -3.159495e-11, 5.08209e-11, 8.099099e-11, 
    -2.527245e-11, -9.136714e-11, -1.199019e-11, -8.429035e-12, 
    -4.476131e-11, 1.010969e-12, -2.382716e-12, -2.287281e-12, -2.94742e-12, 
    2.756684e-12, 9.581891e-12, 5.10858e-12, 3.758216e-11, -1.480793e-11, 
    7.216161e-11, -6.62026e-12, -8.882894e-12, -1.387801e-11, 5.122347e-12, 
    9.85545e-12, 4.532441e-11, -5.204059e-12, -5.632161e-12, 2.911227e-12, 
    3.394396e-12, 1.220652e-10, -3.460343e-12, 1.675882e-13, -3.236988e-11, 
    6.524692e-12, -1.836429e-11, 1.585199e-11, -2.041367e-12, -3.266415e-12, 
    -1.436828e-11, -5.261458e-11, 2.647438e-12, 5.983769e-12, -4.062972e-13, 
    -3.269607e-14, 3.680722e-12, -3.671974e-11, 1.047962e-12, -4.018563e-13, 
    7.140732e-13, -2.153833e-14, 9.39242e-11, 4.290168e-12, -3.284262e-12, 
    3.345424e-11, -1.048428e-11, 3.856693e-12, -1.749911e-11, -3.761658e-12, 
    -3.149436e-12, 2.179175e-10, -8.237566e-11, 5.700351e-11, -3.231482e-11, 
    -8.786971e-12, -8.903389e-11, -1.608291e-11, 3.212786e-11, 1.303913e-11, 
    4.015943e-12, -6.041834e-13, -4.386491e-13, 8.061662e-12, -8.920864e-13, 
    1.472489e-11, 1.307399e-12, 7.88554e-11, 2.979839e-13, 5.3898e-11, 
    -2.747114e-11, 4.53475e-11, 2.054468e-11, -4.430012e-12, 2.044892e-14, 
    7.798207e-13, 7.159828e-12, -2.308078e-11, -2.198353e-12, -2.590017e-12, 
    -1.121812e-10, 2.345679e-13, 6.24878e-13, 3.214096e-12, -1.75191e-11, 
    -4.742829e-12, -1.276868e-11, -3.153319e-11, 2.096268e-12, 1.35586e-13, 
    -3.991496e-11, -1.422884e-11, -9.041878e-12, 3.680678e-11, 1.914624e-11, 
    1.20195e-11, -2.289946e-12, -8.057999e-13, 2.706724e-13, 5.13567e-12, 
    1.112199e-11, -3.366196e-14, 2.822187e-13, 2.346179e-13, 1.240347e-11, 
    6.950218e-12,
  9.585888e-12, -3.618106e-11, 5.297429e-11, 1.564333e-10, 1.867633e-10, 
    9.211187e-11, -1.469691e-11, -8.412671e-11, 8.091283e-11, 4.219134e-10, 
    -2.136973e-10, -5.325185e-11, 3.073919e-11, -2.743916e-11, -7.229439e-11, 
    2.09166e-13, -1.942135e-12, -4.575229e-12, -6.481038e-12, -9.890533e-12, 
    -6.538103e-12, 1.350942e-11, 1.397482e-11, -5.812262e-11, 2.18503e-11, 
    6.62006e-11, -3.217582e-11, -3.562861e-11, 2.049316e-11, 4.333267e-11, 
    6.000511e-11, 7.286549e-11, -1.006317e-10, 3.29814e-11, 7.374346e-11, 
    1.260532e-10, -2.391065e-12, -3.869127e-14, -6.922618e-11, 4.489476e-12, 
    -2.74174e-11, 1.282507e-11, -9.456325e-12, -4.992257e-13, -3.797118e-11, 
    -6.935119e-12, 1.411538e-12, 5.884071e-12, -5.81184e-12, -2.158829e-13, 
    7.945367e-12, -3.728196e-11, 2.492096e-12, 9.228618e-13, 1.29563e-13, 
    4.449774e-13, -3.265366e-11, 7.5282e-13, 2.279243e-12, 2.525258e-12, 
    -9.41891e-12, 1.430878e-11, -4.943135e-11, -5.272183e-12, -3.736167e-12, 
    1.816096e-10, -4.254692e-10, 1.517366e-10, -1.095344e-10, -3.348455e-11, 
    -1.44744e-10, -4.158296e-11, -8.437007e-11, -1.264122e-11, -4.895506e-12, 
    1.396661e-13, -1.466605e-13, 6.933232e-12, -1.909561e-12, 2.418932e-11, 
    -2.772227e-12, 1.239608e-10, -1.379341e-12, 6.765322e-11, -2.249956e-11, 
    1.098408e-10, 9.375833e-12, 7.716272e-12, 1.826386e-13, 4.369838e-13, 
    -1.13356e-11, -1.918266e-11, -2.135958e-12, -2.755667e-11, -1.644997e-10, 
    7.650503e-12, 3.21978e-12, 2.784639e-11, -1.098122e-11, -4.259304e-12, 
    -5.833334e-12, -1.170142e-11, 3.403389e-12, -4.575229e-13, -6.982348e-11, 
    -1.503575e-11, 4.509126e-11, 6.923151e-11, 1.051226e-11, 1.229616e-11, 
    2.905898e-12, 8.667067e-12, -4.719558e-12, -6.405987e-13, 3.774914e-11, 
    7.398527e-14, -3.431699e-13, 6.556561e-13, 6.28031e-12, 1.65683e-11,
  -4.333844e-11, -1.528044e-11, 1.023188e-10, 1.62274e-10, 1.047324e-10, 
    -1.782774e-11, -6.726819e-11, 1.226745e-10, 2.508582e-10, 2.62337e-10, 
    -2.193474e-10, -2.281442e-11, 9.64806e-12, -1.244029e-10, -2.022194e-10, 
    3.974598e-14, -1.66529e-12, -9.505063e-12, -1.134809e-11, -6.186385e-12, 
    7.060352e-12, 1.084843e-11, -7.510814e-11, -2.360443e-10, -4.628409e-11, 
    1.991596e-10, 4.077116e-11, -7.678502e-11, 8.10465e-11, 1.096903e-10, 
    4.633294e-11, 8.739742e-11, -4.289258e-11, 6.295653e-11, 5.92193e-13, 
    3.392644e-10, 2.094991e-12, -4.141132e-14, -2.559888e-10, -6.898038e-13, 
    -2.592002e-11, 5.957235e-12, -4.544698e-12, 2.556955e-12, -5.307998e-11, 
    -3.244316e-11, 1.159739e-12, -6.478151e-13, -2.237868e-11, 9.769685e-13, 
    1.723577e-11, -4.645062e-11, 2.859935e-14, -1.105738e-12, -2.664535e-15, 
    1.982858e-13, -7.064904e-11, -4.017675e-13, 4.6529e-12, 6.343237e-11, 
    -3.143197e-11, 2.274958e-11, -7.497047e-11, -7.547163e-12, -5.199263e-12, 
    1.486649e-10, 1.816722e-10, 4.635534e-10, -4.481326e-11, -8.372036e-11, 
    -1.18068e-10, 8.135936e-12, 2.223455e-10, -8.265233e-11, -1.353739e-11, 
    6.32161e-13, -7.549517e-15, 1.330092e-11, -1.850808e-12, 2.940692e-11, 
    -5.622169e-12, 1.073157e-10, -3.628653e-12, 6.453926e-11, -1.00544e-11, 
    2.224188e-10, 2.813727e-11, 1.333489e-11, -3.736803e-13, 9.383605e-13, 
    -4.086975e-11, -8.728618e-12, -1.441069e-12, -2.977165e-11, 
    -1.705052e-10, 7.088819e-12, 1.170082e-11, 2.518097e-11, -1.248224e-11, 
    -4.629941e-12, -9.233725e-12, 1.284917e-12, 4.059808e-12, 1.523226e-13, 
    -3.778422e-11, 1.874279e-12, 1.281346e-10, 4.78344e-11, -1.377676e-11, 
    1.141198e-11, 2.167821e-12, 2.285883e-11, -1.066147e-11, 1.075606e-11, 
    7.786594e-11, 1.314504e-13, -1.081468e-12, 5.800915e-14, 3.309825e-12, 
    4.364487e-11,
  -6.611023e-11, -1.105338e-12, 8.745937e-11, 1.303904e-10, -2.305267e-12, 
    -9.306289e-11, -1.522293e-11, 5.306142e-10, 3.186353e-10, -2.782818e-10, 
    -1.046314e-10, -1.031704e-10, -4.453105e-11, -2.221872e-10, -3.82316e-10, 
    -7.626788e-13, -1.915179e-12, -9.706902e-12, -1.152667e-11, 6.146639e-12, 
    3.481704e-11, 8.255618e-13, -7.266765e-11, -3.636775e-10, -6.046319e-11, 
    1.584488e-10, 3.044232e-12, -7.094014e-11, 6.205125e-11, 1.814038e-10, 
    1.223674e-10, -3.628786e-11, 1.269718e-10, 1.244467e-10, -6.953993e-12, 
    1.343001e-10, 6.384226e-12, 1.088019e-14, -5.734857e-10, -7.909851e-12, 
    -1.354001e-11, -8.032242e-12, 7.987611e-12, -1.051798e-13, -2.205653e-10, 
    -8.378231e-11, -4.43201e-13, -9.788392e-12, -5.789884e-11, 4.666989e-12, 
    1.808731e-11, -9.040724e-11, -1.171596e-12, -9.540192e-12, -9.232614e-14, 
    -3.703704e-13, -1.370712e-10, -5.536017e-13, -1.119025e-11, 1.685951e-10, 
    -6.604362e-11, 2.939649e-11, -4.190204e-11, -6.775469e-12, -5.045831e-12, 
    1.658411e-10, 6.845502e-11, 6.656999e-10, -3.945066e-11, -1.059344e-10, 
    -4.623368e-11, 3.368461e-11, 1.76946e-10, -1.096736e-10, -3.241496e-12, 
    2.811085e-13, 1.600942e-13, 2.149836e-11, 1.558997e-12, 2.618661e-11, 
    -7.904788e-12, 8.499196e-11, -4.177991e-12, 1.006439e-11, 1.577605e-10, 
    2.823666e-10, -1.122396e-10, 2.275646e-11, -4.449913e-13, 3.33733e-12, 
    -5.169776e-11, -8.303669e-12, -7.085443e-13, -1.104032e-11, 
    -1.257248e-10, 4.70557e-13, 2.376792e-11, 1.089577e-10, -3.784129e-11, 
    -5.775913e-12, -1.107692e-11, 2.03112e-11, 2.908729e-12, 2.11392e-12, 
    -3.262413e-11, 1.875256e-11, 1.078457e-10, -7.177325e-11, -3.489697e-11, 
    1.036637e-11, 1.883382e-12, 3.455591e-11, 2.831957e-12, 2.504352e-11, 
    1.138507e-10, 5.035972e-14, -5.898615e-13, -7.011058e-14, 2.550626e-12, 
    8.982903e-11,
  -6.185541e-11, -3.45981e-11, 7.606715e-11, 9.795631e-11, -7.125855e-11, 
    -5.047163e-11, 1.028662e-10, 8.241434e-10, 5.375966e-10, -1.594893e-10, 
    -5.427658e-11, -3.503127e-10, 4.862866e-11, -3.079892e-10, -4.073346e-10, 
    -2.739142e-12, -2.301537e-12, -5.46807e-12, 1.774692e-12, 2.70024e-11, 
    4.353229e-11, 8.219203e-12, 1.902221e-10, -3.142766e-10, -9.138823e-11, 
    -4.831779e-11, -1.33296e-10, -2.587441e-11, -5.469225e-11, 2.310747e-10, 
    7.336691e-10, 6.661516e-11, 4.568168e-11, 2.995568e-10, 1.168505e-10, 
    9.2209e-10, 9.203128e-12, -4.32987e-15, -3.363576e-10, -1.447225e-11, 
    4.248157e-12, -4.362644e-11, 1.621236e-11, -1.585204e-12, -3.474909e-10, 
    -2.516209e-11, -6.21192e-12, -1.592748e-11, -9.039507e-11, 6.89071e-12, 
    8.418155e-12, -1.319567e-10, 3.720402e-12, -1.54408e-11, -2.804645e-13, 
    -6.12399e-13, -2.091785e-10, -1.853806e-12, -3.527241e-11, 3.032813e-10, 
    -8.003997e-11, 2.252154e-11, -3.090861e-13, -4.795453e-12, -7.122836e-12, 
    1.360778e-10, 1.776224e-10, 8.747065e-10, -1.900053e-10, -1.532134e-10, 
    -6.538947e-11, 1.114362e-10, -3.826628e-11, -1.082743e-10, 9.494627e-12, 
    -6.026291e-12, 3.612666e-13, 8.240075e-12, 8.154144e-12, 2.724043e-12, 
    -1.126343e-11, 6.690879e-11, -4.764633e-12, -3.317613e-11, 2.824683e-10, 
    2.188525e-10, -4.421503e-10, 1.957456e-11, 2.673917e-12, 1.072209e-11, 
    -1.097584e-10, 3.728466e-11, -4.396483e-14, -1.379448e-11, -2.795897e-11, 
    -8.911095e-13, 4.244427e-11, 2.941647e-10, -6.35092e-11, -8.505908e-12, 
    -6.180745e-11, 5.543294e-11, 4.60576e-13, 4.279799e-12, -1.217249e-10, 
    -1.343281e-11, 1.080025e-12, -1.337135e-10, -2.71756e-11, 1.602363e-11, 
    8.396839e-12, 4.745537e-11, 3.191669e-11, 3.891998e-11, 1.312781e-10, 
    1.483258e-14, 1.158518e-12, 4.145018e-13, 1.838807e-12, 1.197895e-10,
  -4.917311e-11, -7.643308e-11, 8.135714e-11, 9.327827e-11, -2.385292e-11, 
    5.921308e-11, 9.823431e-11, 8.570922e-10, 1.205025e-09, -4.846967e-11, 
    -9.640466e-11, -9.632188e-10, 2.156657e-10, -3.868852e-10, -3.452669e-10, 
    -6.053646e-12, -8.098411e-13, 2.342126e-12, 1.719136e-11, 5.037393e-11, 
    4.271428e-11, 3.496936e-11, 2.840324e-10, 3.368186e-10, -2.886242e-10, 
    -3.156124e-10, -2.388614e-10, -5.850964e-11, -2.050324e-10, 2.575735e-10, 
    1.361578e-11, 2.812399e-10, -3.996821e-10, 4.349658e-10, 1.22057e-10, 
    2.404956e-10, 6.899015e-12, -9.392487e-14, 1.987388e-11, -1.73511e-11, 
    -5.48301e-11, -1.401794e-10, 2.408296e-11, -1.223716e-12, -6.217054e-10, 
    3.010037e-11, -2.26823e-11, -1.803802e-11, -1.004356e-10, 1.618816e-12, 
    2.224221e-12, -6.557244e-11, 5.333867e-12, -8.592593e-12, -1.753264e-13, 
    -1.262102e-12, -4.809966e-10, -9.049472e-12, -6.366196e-11, 2.608362e-10, 
    -8.490453e-11, -1.92717e-11, 8.381029e-11, -6.788525e-12, -1.624087e-11, 
    3.356604e-11, -1.153252e-09, 2.525027e-09, -4.351595e-10, -2.225562e-10, 
    -2.081091e-10, 3.30969e-10, -5.683152e-10, -6.144596e-11, 9.760193e-12, 
    -1.799272e-11, 3.601563e-13, -3.467981e-11, 2.218425e-11, 1.491962e-11, 
    -1.792788e-11, 2.735354e-11, -7.841727e-12, -6.810019e-11, 5.060752e-10, 
    1.555733e-10, -5.260681e-10, 3.542056e-12, 1.351919e-11, 2.784528e-11, 
    -2.619576e-10, 1.415401e-10, 1.414868e-12, -6.152074e-11, -1.310738e-10, 
    -3.631282e-11, 7.292798e-11, 3.909193e-10, -6.971135e-11, -3.605649e-12, 
    -7.73035e-11, 1.496953e-10, -2.259082e-12, 4.026224e-12, -2.704894e-10, 
    -1.962785e-10, -1.567049e-10, 2.118892e-10, 3.315215e-11, 1.868905e-11, 
    7.313261e-12, 8.028067e-11, 5.859491e-11, 4.996714e-11, 1.167635e-10, 
    3.678835e-13, 3.461675e-12, 2.10304e-12, -6.724621e-13, 1.174438e-10,
  -3.668532e-11, -7.963763e-11, 1.327987e-10, 2.414833e-10, 1.564011e-10, 
    8.889423e-11, -3.853096e-11, 3.855813e-10, 1.567388e-09, 9.809824e-10, 
    -1.589537e-10, -1.00102e-09, 3.202238e-11, -4.61684e-10, -4.803642e-10, 
    -7.874768e-12, 2.938449e-12, 1.845013e-11, 2.592504e-11, 6.57181e-11, 
    4.431833e-11, 5.840661e-11, 2.145804e-10, 1.163469e-09, -6.831513e-10, 
    -4.867005e-10, -3.319354e-10, -3.454961e-10, -7.283383e-10, 2.887699e-10, 
    -1.497469e-10, 2.210214e-10, -9.85537e-10, 8.577175e-10, 1.038103e-10, 
    1.904324e-09, 1.860929e-11, -3.175238e-14, 1.295923e-10, -1.698517e-11, 
    2.094154e-10, -2.611191e-10, 3.949063e-11, -2.462058e-12, -7.947811e-10, 
    3.012577e-10, -5.251977e-11, -2.086775e-11, -8.36625e-11, -1.476352e-11, 
    4.374723e-12, 9.731771e-11, -1.109601e-11, 8.067147e-12, -7.490453e-13, 
    -2.845724e-12, -6.427623e-10, -2.784013e-11, -2.390348e-10, 2.282781e-10, 
    -8.858336e-11, -9.482903e-11, 1.991918e-10, -1.286544e-11, -2.495106e-11, 
    -1.278e-10, -6.327614e-10, 3.87128e-09, -9.867449e-10, -4.251763e-10, 
    -1.909832e-10, 4.449312e-10, -2.026557e-10, -9.507062e-12, 7.883471e-13, 
    -3.059952e-11, 4.474199e-13, -9.557244e-11, 4.223644e-11, 1.377565e-11, 
    -3.24345e-11, -1.080278e-11, -1.230038e-11, -1.455476e-10, -9.341861e-11, 
    -1.080274e-10, 6.911449e-11, -9.903189e-12, 3.467213e-11, 5.002754e-11, 
    -5.033129e-10, -1.450527e-10, 4.547918e-12, -7.694644e-12, -1.825633e-10, 
    -1.273554e-10, 1.138329e-10, 4.804761e-10, -5.934808e-11, 2.843237e-12, 
    7.405099e-11, 3.031184e-10, -6.254108e-12, 1.552314e-12, -3.362697e-10, 
    -4.414442e-10, -4.05544e-10, 8.117205e-10, 1.833378e-10, -3.42304e-12, 
    8.331114e-12, 1.135092e-10, 8.089884e-11, 3.56728e-11, 7.335998e-11, 
    2.216005e-12, 5.715428e-12, 5.149825e-12, -5.651368e-12, 8.425083e-11,
  -1.478284e-11, -1.417995e-10, 2.336229e-10, 5.068017e-10, 3.629275e-10, 
    2.085336e-10, -5.529799e-11, -2.227161e-10, -1.270735e-10, 2.108731e-09, 
    -1.384599e-10, 8.956391e-11, -1.006907e-09, -5.036647e-10, -5.664731e-10, 
    2.438583e-12, 5.74687e-12, 4.775202e-11, 2.605027e-11, 7.248957e-11, 
    4.91589e-11, 3.41096e-11, 2.453966e-10, 1.362803e-09, -5.548699e-10, 
    -5.034302e-10, -2.968612e-10, 2.268798e-10, -1.095831e-09, 3.048726e-10, 
    3.647571e-11, -2.315907e-10, -1.72161e-10, 1.827992e-09, 2.628653e-11, 
    3.600736e-09, 1.857394e-11, 5.622169e-13, -7.539569e-11, -1.517968e-11, 
    -6.323831e-12, -2.867786e-10, 5.750422e-11, -1.148343e-11, -1.112518e-09, 
    1.371507e-09, -7.926459e-11, -2.602452e-11, -7.158789e-11, -1.996869e-11, 
    -9.204282e-11, 3.757066e-10, -1.871179e-11, 4.775487e-11, 5.595524e-14, 
    -4.126477e-12, 4.670504e-10, -6.753211e-11, -8.310142e-10, 3.326273e-11, 
    -3.871747e-11, -1.705018e-10, 2.301235e-10, -8.319035e-12, -2.664464e-11, 
    -2.474749e-10, -1.272245e-09, -3.290523e-10, -1.909356e-09, 
    -7.872138e-10, 4.317791e-10, 8.136745e-10, -1.468408e-09, -5.784884e-11, 
    -1.799876e-11, -3.754508e-11, 7.96252e-13, -1.450315e-10, 5.666747e-11, 
    -2.655227e-10, -5.987388e-11, -3.924585e-11, -1.818456e-11, 4.064766e-10, 
    -5.049614e-10, -7.691661e-10, 1.413373e-09, -1.899991e-11, 5.372514e-11, 
    7.184831e-11, -9.119852e-10, -4.558998e-10, 7.896794e-12, 2.697469e-10, 
    -3.887912e-10, -2.237268e-10, 1.668759e-10, 5.71287e-10, -3.079137e-11, 
    -6.495071e-12, 2.000924e-10, 5.201122e-10, -1.11795e-11, 4.766187e-12, 
    -2.178773e-10, -5.325269e-10, -6.642544e-10, 8.610073e-10, 4.843947e-10, 
    -1.022649e-10, -1.804068e-11, 1.060805e-10, 1.230553e-10, 7.442935e-11, 
    2.798828e-11, 5.056222e-12, 1.027312e-11, 8.185674e-12, -7.559731e-12, 
    2.413358e-11,
  3.891643e-11, -2.758398e-10, -2.065619e-10, 4.607443e-10, 4.805116e-10, 
    3.92042e-10, 2.765077e-10, -3.433414e-10, -8.83837e-10, 1.585008e-09, 
    -6.31843e-10, 2.332925e-10, -6.319425e-10, -4.976428e-10, -6.870309e-10, 
    3.351631e-12, -1.509193e-11, 8.099477e-11, 6.843415e-12, 9.253398e-11, 
    6.185275e-11, -5.81224e-12, 2.903491e-10, 1.309999e-09, -7.206111e-10, 
    -3.503686e-11, -9.243735e-10, 5.716956e-10, -4.759286e-10, 3.996234e-10, 
    -1.016247e-09, -4.122356e-10, -3.251586e-10, 3.223683e-09, 1.331841e-10, 
    6.03594e-09, 2.753211e-11, 1.522338e-12, -1.495835e-10, -2.90612e-12, 
    -6.1398e-11, -2.114788e-10, 4.076028e-11, -6.397205e-11, -1.458588e-09, 
    2.139977e-09, -6.202683e-11, -2.691181e-11, -1.417504e-10, -2.097877e-12, 
    -3.848957e-10, 3.760974e-10, -4.390159e-11, 1.151733e-10, 1.297735e-11, 
    -2.316369e-12, 1.619924e-09, -1.405638e-10, -1.980833e-09, -2.097931e-10, 
    2.223999e-12, -2.357794e-10, 6.100009e-11, 2.774669e-11, -8.439826e-12, 
    -3.490257e-10, -5.294325e-10, 2.062066e-10, -1.917421e-09, -1.081972e-09, 
    1.182791e-09, 1.641276e-09, 4.838796e-11, -4.328697e-10, -6.261232e-11, 
    -3.020517e-11, 1.517009e-12, -1.590763e-10, 3.454854e-11, -9.402541e-10, 
    -1.016573e-10, -2.263345e-11, -3.165468e-11, 8.592238e-10, -5.604832e-10, 
    -7.391918e-10, 2.715765e-09, -2.855671e-11, 6.215661e-11, 3.003464e-10, 
    -1.337455e-09, -4.239226e-10, 5.25624e-12, 5.64787e-10, -1.144286e-09, 
    -2.828642e-10, 2.652058e-10, 6.285887e-10, -3.007727e-11, -2.727489e-11, 
    1.146816e-11, 7.002705e-10, -1.036105e-11, 2.209388e-11, 1.148095e-10, 
    -4.449632e-10, -5.234995e-10, 1.222062e-09, 1.403095e-09, 6.524914e-11, 
    -9.528378e-11, -1.028155e-11, 2.011546e-10, 1.284874e-10, -3.444001e-11, 
    7.425172e-12, 1.703615e-11, 9.823919e-12, -9.225065e-12, -4.635581e-11,
  -9.627854e-13, -1.912888e-10, -1.92923e-10, 9.487913e-10, 1.354334e-09, 
    4.584244e-10, 5.815046e-10, -3.243379e-10, -3.907381e-10, -1.694112e-10, 
    -1.167574e-09, 2.520117e-10, -1.829942e-09, -4.464162e-10, -6.191208e-10, 
    -1.737063e-11, -2.870053e-10, 9.101697e-11, -1.99547e-11, 1.232117e-10, 
    9.398704e-11, 1.514522e-11, 2.468674e-10, 9.19389e-10, -3.709236e-09, 
    1.653039e-09, -1.531735e-09, -8.179804e-10, 5.752732e-10, 1.286768e-09, 
    3.781285e-09, -1.860133e-09, -6.309655e-10, 4.153893e-09, -1.050431e-10, 
    4.884338e-09, -1.146674e-11, 3.572254e-12, -1.006306e-10, -1.953353e-11, 
    3.569838e-11, -1.897611e-10, -1.069544e-11, -2.636422e-10, -1.781093e-09, 
    1.518213e-09, -4.138911e-12, -9.202417e-11, -3.33096e-10, 6.58269e-11, 
    -5.762022e-10, -4.10477e-10, -7.609842e-11, 1.899316e-10, 2.897647e-11, 
    4.828138e-12, 2.703228e-09, -2.475318e-10, -3.421808e-09, -3.243557e-10, 
    3.431566e-11, -2.909211e-10, -2.603784e-11, 6.489742e-11, 2.467786e-11, 
    -4.479368e-10, 4.322764e-10, 3.873275e-10, -7.472174e-10, -1.559425e-09, 
    8.012968e-10, 2.046679e-09, 2.396838e-10, -9.85704e-10, -1.536762e-10, 
    -1.535128e-11, 5.15854e-12, -1.478337e-10, -1.194262e-11, -7.064571e-11, 
    -1.193072e-10, 1.845382e-10, -5.691803e-11, 1.928381e-09, 8.036967e-09, 
    1.068468e-09, 3.202882e-09, -1.635314e-11, 1.362205e-10, 1.052815e-09, 
    -2.240423e-09, -1.286701e-10, -1.630696e-12, 1.792081e-10, 1.021156e-10, 
    -3.928946e-10, 4.015512e-10, 9.100098e-10, -1.383818e-10, -5.456045e-11, 
    -7.903012e-11, 7.864789e-10, -2.073008e-12, 5.508172e-11, 2.18332e-10, 
    -1.457074e-10, -1.482157e-10, 6.396483e-10, 1.354028e-09, 8.395951e-10, 
    -1.261249e-10, -2.755023e-10, 2.282299e-10, 2.155964e-10, -1.066702e-10, 
    1.324665e-11, 2.514255e-11, 1.193778e-11, -8.230305e-12, -1.134559e-10,
  1.542766e-10, -8.779111e-11, 3.580642e-09, 1.491419e-09, 2.816055e-09, 
    1.21641e-09, 4.379537e-10, 2.266809e-10, -6.665957e-11, -1.652065e-09, 
    -8.576073e-10, 5.228529e-11, -3.441965e-09, -3.174527e-10, -3.319904e-10, 
    -4.292178e-11, -6.463886e-10, 6.056311e-11, -2.925127e-11, 1.342251e-10, 
    1.532676e-10, 8.641976e-11, 1.978044e-10, 8.769412e-10, 1.071676e-10, 
    3.435677e-09, -4.613945e-10, 1.421263e-10, -4.019647e-10, 2.163578e-09, 
    4.824106e-09, -1.288894e-08, -1.090424e-09, 3.626841e-09, -3.034692e-10, 
    2.762835e-09, -1.32048e-10, 2.000178e-12, 1.538076e-10, -2.768935e-10, 
    6.772964e-11, -3.30683e-10, -4.093792e-11, -4.061909e-10, -2.157545e-09, 
    4.217249e-10, 1.013589e-11, -4.45997e-10, -4.683663e-10, 2.102887e-10, 
    3.872103e-11, -6.900329e-10, 6.841605e-11, 2.238586e-10, 2.288942e-11, 
    1.65663e-11, 1.226116e-09, -3.838245e-10, -4.682644e-09, 1.264731e-10, 
    2.984635e-11, -3.204939e-10, -8.700951e-11, -1.074618e-10, 3.271125e-11, 
    -6.110064e-10, 4.145608e-09, -3.682707e-10, 1.96426e-10, -2.277002e-09, 
    -9.156729e-10, 1.306123e-09, 3.387619e-10, -8.803163e-10, -1.476785e-10, 
    -1.295675e-11, 9.972467e-12, -1.291518e-10, -4.660663e-11, 4.473186e-10, 
    -5.254819e-11, 5.678043e-10, -8.761347e-11, 3.253479e-09, 4.281564e-09, 
    1.197808e-09, 2.485368e-09, -2.810197e-12, 4.642049e-10, 2.064159e-09, 
    -1.711211e-09, -3.476792e-10, -6.06093e-12, -4.268779e-09, 1.023327e-09, 
    -6.928325e-10, 4.933532e-10, 1.448303e-09, -3.370495e-10, 3.769429e-12, 
    -6.773959e-11, 7.7205e-10, -1.027001e-11, 8.751666e-11, -4.639098e-10, 
    -3.333831e-10, 2.976073e-10, 6.584351e-10, 6.895e-10, 2.324175e-09, 
    -2.846079e-11, -5.393836e-10, -5.419665e-11, -6.536247e-10, 
    -2.919727e-10, 2.140084e-11, 3.3058e-11, 2.229861e-11, -6.442846e-12, 
    -1.785843e-10,
  3.440341e-10, 2.009774e-09, 3.43551e-10, -5.930438e-10, -2.165319e-09, 
    -1.301355e-09, -1.177593e-09, 1.158316e-09, -6.972662e-10, -1.626045e-09, 
    -6.954046e-10, 9.04226e-10, -1.658517e-09, 1.424674e-10, -8.379537e-10, 
    1.760603e-10, -3.371859e-10, -2.84718e-10, -4.037659e-12, 1.433769e-10, 
    2.587548e-10, 2.163496e-10, 1.721823e-10, 1.414353e-09, 4.772208e-09, 
    3.610911e-09, 1.831427e-09, 2.309083e-09, -4.991101e-10, -3.932854e-12, 
    6.23459e-09, -1.720641e-08, -1.257305e-11, 1.39406e-09, -7.702532e-10, 
    6.2136e-09, -2.615202e-10, 3.751666e-12, -4.185733e-09, -1.014265e-09, 
    3.933344e-10, -6.407639e-10, -1.415401e-11, -1.955671e-10, -2.372428e-09, 
    -3.616627e-10, -1.596696e-10, -1.169067e-09, 1.434799e-11, 1.239568e-10, 
    6.261995e-10, -6.598349e-10, -1.781542e-11, 2.215991e-10, -7.822365e-12, 
    2.144063e-11, -8.579768e-10, -5.546404e-10, -4.609259e-09, -2.743175e-09, 
    2.238565e-11, -3.466134e-10, -3.595737e-10, -1.038861e-09, -1.578506e-10, 
    -3.838743e-10, 5.642637e-09, -3.433893e-09, -9.972823e-11, -2.578314e-09, 
    -2.377913e-09, 2.044978e-10, 3.373266e-10, 7.579537e-10, 1.420396e-10, 
    -2.355804e-11, 7.574386e-12, -1.510685e-10, -1.679975e-10, -3.815259e-11, 
    8.35918e-11, 1.014278e-09, -1.171792e-10, 5.331717e-09, 3.095455e-09, 
    2.304184e-10, 9.536798e-10, 8.629542e-12, 1.535907e-09, 2.51649e-09, 
    -2.326139e-10, -1.18081e-09, -4.323653e-12, -9.223756e-09, 1.606114e-09, 
    -1.110106e-09, 4.801912e-10, 2.479798e-09, -4.689262e-10, -1.77117e-11, 
    -8.551773e-10, 5.585434e-10, -5.399237e-11, 9.83551e-11, 2.579625e-11, 
    5.789396e-10, -2.487965e-11, -2.921716e-10, 9.521877e-10, 4.830074e-09, 
    2.846043e-10, -6.178418e-10, -2.220979e-10, 3.96529e-10, -6.065299e-10, 
    3.083258e-11, 3.69873e-11, 4.67022e-11, -8.592238e-12, -2.382556e-10,
  1.864535e-10, 7.134453e-09, 9.536002e-09, 5.39476e-09, -1.668533e-08, 
    -7.713872e-09, -5.06531e-09, 4.250253e-10, 6.091483e-11, -8.072263e-10, 
    -4.309229e-10, 2.337039e-09, -1.903707e-09, 4.488498e-11, -9.815366e-10, 
    -3.824239e-10, 2.374883e-09, -1.350507e-09, 1.391598e-11, 2.31708e-11, 
    2.570815e-10, 4.564029e-10, 1.448726e-10, 1.229218e-09, 5.840839e-09, 
    2.087837e-09, 4.052659e-09, 8.894695e-09, -1.230283e-09, -6.567682e-09, 
    1.476108e-08, -9.045259e-09, -9.588774e-11, -5.518288e-10, -1.57916e-09, 
    9.625303e-09, -3.363382e-10, 7.048584e-12, -1.889184e-09, -1.995188e-09, 
    5.610857e-10, -1.15778e-09, 3.607497e-10, -3.199725e-10, -1.772882e-09, 
    3.663914e-10, -7.728218e-10, -1.850125e-09, 1.153917e-09, 1.289138e-10, 
    1.422958e-09, -2.823342e-10, -1.776996e-10, 2.168477e-10, -3.992966e-11, 
    -7.808865e-12, -2.988251e-09, -7.92177e-10, -4.894274e-09, 7.144301e-09, 
    3.445422e-11, -4.854925e-10, -8.203287e-10, -2.762577e-09, -1.76958e-09, 
    -3.445209e-10, 8.758789e-10, -6.598235e-09, -2.113545e-09, -2.883034e-09, 
    -2.044168e-09, 1.871356e-10, -1.74466e-09, -8.877166e-10, 2.988443e-10, 
    -3.801404e-12, 8.821388e-12, -1.86354e-10, -3.439382e-10, -1.371845e-10, 
    4.125056e-10, 1.6932e-09, -1.257447e-10, 7.178279e-09, 1.68874e-09, 
    6.719247e-10, -1.14246e-09, 1.708855e-11, 3.304476e-09, 3.780862e-09, 
    4.305186e-09, -7.612855e-10, -2.163603e-11, -1.133583e-08, 5.648104e-11, 
    -1.508774e-09, 3.134986e-10, 4.039101e-09, -4.342482e-10, -7.02343e-11, 
    -3.858865e-09, 3.4637e-10, -1.583551e-10, 8.309442e-11, 8.402097e-10, 
    2.602363e-10, -2.061071e-10, 1.164103e-09, 2.219089e-09, 7.148778e-09, 
    1.660183e-10, -5.562057e-10, -2.517524e-10, 9.05608e-10, -9.842935e-10, 
    4.480825e-11, 3.931078e-11, 7.968293e-11, -4.339817e-11, -3.403429e-10,
  -2.519585e-10, 1.06273e-08, 1.012009e-08, 8.805443e-09, 4.292446e-09, 
    2.473087e-09, -6.837297e-09, -3.435645e-09, 2.06478e-09, -2.070806e-10, 
    7.417782e-10, -1.181263e-09, -2.358689e-09, 9.452776e-10, -1.302794e-09, 
    -8.040644e-10, 5.248444e-09, -1.276561e-09, 1.110578e-11, -2.031868e-10, 
    2.960121e-10, 8.151062e-10, 6.804157e-11, 6.853043e-10, 1.758053e-09, 
    -7.274252e-10, 2.059011e-09, 4.32492e-08, 4.574957e-09, -1.310664e-08, 
    2.463446e-08, 5.0361e-09, 1.541281e-09, 1.000274e-09, -1.850992e-09, 
    1.257322e-08, -3.13679e-10, 9.706014e-12, -1.116095e-08, -1.765727e-09, 
    1.517054e-09, -1.521045e-09, 4.081571e-10, -5.068985e-10, -1.040539e-08, 
    -8.384404e-11, -2.211195e-09, -2.056375e-09, 1.795934e-09, 1.167599e-10, 
    2.183629e-09, 2.24162e-10, -6.611458e-11, 2.762533e-10, -4.209042e-11, 
    -8.35314e-11, -5.879428e-09, -1.154703e-09, -6.765663e-09, 9.650957e-09, 
    -3.66839e-10, -8.125198e-10, -9.837322e-10, -3.660307e-09, -7.553155e-09, 
    5.112696e-09, 3.65398e-09, -5.201429e-09, 1.649141e-09, -8.451195e-10, 
    -2.210186e-09, 7.950121e-10, -6.469719e-09, -4.493074e-09, 5.010435e-10, 
    5.010747e-11, 1.638512e-11, -1.873275e-10, -4.289483e-10, 7.866277e-10, 
    9.067378e-10, 2.590755e-09, -1.453913e-10, 8.11653e-09, -2.956682e-09, 
    1.810548e-09, -5.625537e-09, 8.91589e-11, 5.25816e-09, 5.049628e-09, 
    1.180496e-08, -3.182663e-10, -4.436629e-11, -5.905095e-09, -2.996757e-09, 
    -2.751005e-09, 2.062961e-10, 4.871168e-09, -3.11843e-10, -5.716742e-11, 
    -4.530534e-09, 2.675122e-10, -3.821334e-10, 5.761081e-11, 7.266294e-10, 
    5.761081e-10, 1.440327e-09, 3.943939e-09, 9.905534e-10, 6.895476e-09, 
    3.432774e-10, -5.239542e-10, -4.679919e-10, 1.281819e-10, -1.435183e-09, 
    7.732979e-11, 4.632383e-11, 1.100089e-10, -9.54401e-11, -5.065033e-10,
  -1.035403e-10, 1.007905e-08, 4.139793e-09, 2.177785e-09, 4.572939e-09, 
    2.733486e-09, -4.159489e-09, -1.088722e-08, 9.95442e-10, 1.710134e-10, 
    1.925514e-09, -4.178389e-09, -1.239783e-09, 2.942386e-09, -2.505232e-09, 
    -7.121486e-10, 6.152135e-09, 1.065516e-09, -1.448086e-11, 3.911396e-10, 
    6.3838e-10, 1.263174e-09, 1.132605e-10, 2.498552e-10, 4.206981e-10, 
    2.3025e-09, -3.649603e-09, 3.564324e-08, 9.599177e-09, -1.236566e-08, 
    2.732241e-08, 2.899185e-09, 1.693081e-09, 1.849884e-09, -5.892673e-10, 
    1.703057e-08, -3.390823e-10, 1.661959e-11, -1.133984e-08, -1.348909e-09, 
    4.488106e-09, -1.754614e-09, -1.638014e-10, -7.863554e-10, -1.436163e-08, 
    6.494645e-10, -5.69446e-09, -2.968619e-09, 1.968652e-09, 9.065104e-11, 
    1.775092e-09, 5.93559e-10, 1.479947e-10, 4.283493e-10, -1.864535e-11, 
    -1.431317e-10, -9.34449e-09, -1.67399e-09, -8.780921e-09, 6.727277e-09, 
    -1.064507e-09, -9.227961e-10, -9.377743e-10, -2.680434e-09, 
    -1.155162e-08, 2.570715e-09, 4.850904e-09, -5.024788e-09, 2.167553e-09, 
    1.652069e-09, -6.335767e-10, 8.929248e-10, -4.337068e-09, -3.420837e-10, 
    7.023516e-10, 6.031087e-11, 1.8062e-11, -1.950937e-10, -4.770129e-10, 
    -2.103178e-09, 1.287162e-09, 3.375781e-09, -1.568026e-10, 1.146211e-08, 
    -9.940919e-09, 3.40782e-09, -9.834622e-09, 2.208367e-10, 7.654819e-09, 
    7.244026e-09, 1.29823e-08, -6.954792e-11, 3.107914e-11, -5.709762e-09, 
    3.081198e-10, -6.541422e-09, 6.462699e-10, 3.73322e-09, -3.638831e-10, 
    -5.553602e-11, -1.805461e-09, 2.577867e-10, -7.92344e-10, 5.285727e-11, 
    6.077983e-10, 8.007248e-10, 1.955129e-09, 3.357627e-09, -3.446189e-09, 
    7.64183e-09, 1.393403e-09, -2.465299e-10, -1.281308e-09, -2.837623e-09, 
    -2.024279e-09, 8.99405e-11, 5.561063e-11, 8.024426e-11, -1.175025e-10, 
    -5.820482e-10,
  1.016247e-09, 6.680239e-09, 1.019828e-09, -8.180336e-10, 7.199219e-10, 
    2.247589e-10, 5.141487e-10, -1.404032e-08, -1.516526e-09, 1.57911e-09, 
    1.66915e-09, -3.510593e-09, 3.774403e-10, -6.521077e-10, -9.893597e-10, 
    9.470114e-11, 3.668998e-09, 3.412566e-09, -2.096101e-11, 1.274429e-09, 
    4.869207e-10, 1.452008e-09, 6.09532e-10, 1.929266e-10, -1.644821e-09, 
    6.91773e-09, -3.04675e-09, -1.161544e-08, 6.647213e-09, -2.558693e-09, 
    2.498723e-08, 1.180638e-10, 3.115986e-09, 4.363869e-10, 7.879635e-10, 
    2.235134e-08, -7.660333e-10, 3.03686e-11, -1.024455e-08, -2.356336e-09, 
    7.396477e-09, -1.869125e-09, -1.07903e-09, -8.127898e-10, -2.918455e-09, 
    1.336389e-10, -1.35303e-08, -4.487504e-09, 2.216473e-09, 5.404388e-11, 
    8.886545e-10, 4.774847e-11, 5.506877e-10, 6.957748e-10, -2.465583e-11, 
    -9.742962e-11, -1.686016e-08, -2.361412e-09, -1.409548e-08, 2.083937e-09, 
    -2.007425e-09, -5.639436e-10, -6.630785e-10, -3.564571e-09, 
    -7.224378e-09, 3.15822e-09, 6.269602e-09, -1.220519e-08, -9.017981e-09, 
    4.318395e-09, 7.11907e-10, 7.361223e-11, -1.615604e-09, 6.091227e-09, 
    6.57684e-10, 2.50111e-11, 3.385026e-11, -9.225687e-11, -5.58704e-10, 
    -5.267623e-09, 1.63854e-09, 4.009539e-09, -1.987246e-10, 9.848009e-09, 
    -5.682296e-09, 2.877357e-09, -5.897732e-09, 2.982006e-10, 1.123471e-08, 
    1.060931e-08, 9.58903e-09, -4.345226e-10, 1.416112e-10, -9.887135e-09, 
    1.687113e-09, -7.742802e-09, 1.269427e-10, 9.723635e-10, -3.78293e-10, 
    -6.228902e-11, -5.112497e-10, 1.985647e-10, -1.845962e-09, 1.581952e-10, 
    1.356625e-09, 7.941026e-10, 5.918537e-10, 1.910223e-09, -2.456829e-09, 
    1.358757e-08, 2.785953e-09, 2.369234e-10, -2.371905e-09, -2.638956e-09, 
    -2.073648e-09, 3.320793e-11, 1.05544e-10, 1.267075e-11, -9.336532e-11, 
    -6.291998e-10,
  5.239826e-10, 2.070863e-09, 2.203819e-10, -2.303409e-09, 7.972858e-10, 
    -7.765379e-10, 1.622936e-09, -7.682843e-09, -5.970946e-09, 2.302784e-09, 
    1.760384e-09, -5.884885e-09, 4.927756e-10, -2.995534e-09, -5.07714e-09, 
    8.693126e-10, -1.021476e-09, 4.716242e-09, -9.86482e-10, 1.659203e-09, 
    -4.212097e-10, 1.260219e-09, 1.627939e-09, 2.636398e-10, -4.275762e-10, 
    -5.280754e-11, -2.73161e-09, -1.34832e-08, -4.377512e-09, 4.127003e-09, 
    2.719662e-08, -3.021398e-09, 4.90536e-09, -1.185072e-09, -3.690275e-10, 
    2.497046e-08, -1.629314e-09, 6.304646e-11, -1.674113e-08, -3.835032e-09, 
    6.254493e-09, -7.001972e-10, -1.793012e-09, -1.317181e-09, -4.304752e-10, 
    -7.368044e-10, -2.49413e-08, -7.041535e-09, 2.192837e-09, 6.450662e-11, 
    -7.783783e-10, -1.184731e-09, 1.477258e-09, 1.157105e-09, -8.064234e-11, 
    2.55227e-11, -2.869962e-08, -3.867399e-09, -2.69492e-08, -4.19594e-09, 
    -2.323361e-09, -5.352945e-10, -2.524416e-10, -9.273606e-09, 
    -1.567048e-09, 5.316906e-09, 8.97785e-09, -2.250107e-08, -4.589651e-09, 
    1.160004e-09, 1.385843e-09, 1.342812e-09, 4.143317e-10, 5.130062e-09, 
    2.683749e-10, 2.12026e-11, 6.685497e-11, 2.941647e-11, -7.249341e-10, 
    -1.841158e-09, 2.176222e-09, 4.500089e-09, -2.596892e-10, 4.980848e-09, 
    2.251511e-09, 1.525393e-09, 3.551747e-09, 4.417871e-10, 1.610292e-08, 
    1.544763e-08, 8.155723e-09, -9.071641e-10, 2.57856e-10, -7.973309e-09, 
    1.452406e-09, 4.381252e-09, 1.332853e-09, 3.134858e-09, -2.042384e-10, 
    -6.000391e-11, -7.610765e-10, 1.250555e-10, -3.723517e-09, 5.14838e-10, 
    4.595165e-09, -3.115019e-10, 5.574066e-10, -1.209287e-09, -3.444939e-09, 
    1.538189e-08, 1.813589e-09, -9.401901e-11, -2.116678e-09, -5.89597e-09, 
    -1.571834e-09, -3.591935e-11, 2.769056e-10, -9.242029e-11, -5.32836e-11, 
    -5.808829e-10,
  -4.117737e-10, -5.88642e-09, -1.293756e-09, -1.241062e-09, 1.776073e-09, 
    -3.096261e-10, -1.066439e-09, 3.911396e-10, -1.139438e-08, 7.170229e-10, 
    2.044999e-09, -7.359631e-09, -1.084913e-09, -7.059953e-10, -1.221764e-08, 
    -6.540177e-10, -4.069506e-09, 5.277371e-09, -3.600768e-09, 1.165461e-09, 
    -1.173646e-09, 1.304443e-09, 2.577622e-09, 8.124061e-10, -2.197567e-10, 
    -1.850822e-10, 1.433961e-08, -1.042781e-08, -1.002695e-08, 4.609319e-09, 
    2.877289e-08, -4.495234e-09, 7.460187e-09, -4.344599e-09, -9.946007e-09, 
    3.052003e-08, -1.666467e-09, 1.123581e-10, -2.384525e-09, -5.771733e-09, 
    2.576996e-09, 1.816261e-09, -2.222933e-09, -2.017959e-09, -3.431353e-09, 
    -6.772325e-09, -2.648855e-08, -1.061743e-08, 1.250214e-09, 3.002398e-11, 
    -3.512874e-09, -1.707065e-09, 2.592236e-09, 1.837441e-09, 1.253554e-10, 
    9.512746e-11, -3.964328e-08, -3.7939e-09, -3.974915e-08, -1.503749e-08, 
    3.626155e-09, -1.047056e-10, -8.266738e-10, -1.900621e-08, 2.939385e-09, 
    2.914874e-09, 1.374349e-08, -2.986445e-08, -3.002924e-09, -7.143115e-09, 
    5.232437e-10, 7.558754e-09, 1.202807e-09, 2.507136e-09, -3.106038e-10, 
    9.509904e-11, 4.715872e-11, 7.9595e-11, -9.734749e-10, 4.507683e-11, 
    2.708589e-09, 6.354785e-09, -5.20771e-10, -9.208634e-10, 6.591392e-09, 
    1.357989e-09, 4.427477e-09, 8.215579e-10, 1.906178e-08, 2.149864e-08, 
    8.843074e-09, -4.477544e-09, 4.314131e-10, -2.155028e-08, 1.99293e-09, 
    2.62805e-08, 7.031531e-11, 1.360945e-08, 4.053504e-10, -6.144774e-11, 
    -1.819046e-09, -3.816325e-11, -5.264376e-09, 1.078984e-09, 8.633776e-09, 
    -3.16038e-09, 2.501736e-09, -7.435006e-09, 1.950752e-09, 1.263015e-08, 
    1.662215e-09, -1.175295e-09, -3.247465e-09, -1.25267e-08, -4.829474e-09, 
    -4.488925e-11, 5.293828e-10, -1.469083e-10, -3.795719e-11, -4.18197e-10,
  -4.525305e-10, -4.307708e-09, -3.353648e-09, 1.006924e-09, 2.083823e-09, 
    7.369749e-10, -1.931028e-09, 4.810204e-09, -1.354664e-08, -3.896503e-09, 
    2.117304e-09, -6.335654e-09, -2.559034e-09, 4.071978e-09, -2.790784e-09, 
    -2.143361e-09, -5.802798e-09, 4.919087e-09, -6.019071e-09, 3.493597e-10, 
    -4.887966e-10, 1.334968e-09, 2.746674e-09, 1.853039e-09, -6.777441e-10, 
    -7.569838e-10, 2.724164e-09, -9.644509e-09, -8.254347e-09, 1.170298e-08, 
    2.951197e-08, -3.752405e-09, 9.141843e-09, -6.799496e-09, -1.28972e-08, 
    3.689763e-08, -1.853186e-09, 5.501732e-11, -2.231502e-08, -9.672589e-09, 
    -6.616892e-09, 3.670777e-09, -1.785665e-09, -2.575123e-09, -1.123942e-08, 
    -3.624433e-08, -1.947109e-08, -1.353817e-08, -1.755188e-09, 
    -1.565681e-11, -4.704809e-09, -1.642263e-09, 4.561474e-09, 2.819798e-09, 
    7.256119e-10, 1.319904e-10, -4.15406e-08, 1.528917e-10, -2.079796e-08, 
    -2.002157e-08, 7.005838e-09, -3.848868e-10, -2.058073e-09, -2.643999e-08, 
    5.801212e-09, -3.06494e-09, 1.887781e-08, -3.185886e-08, -9.919916e-09, 
    -1.797923e-08, -2.382109e-08, 8.163966e-09, -2.899532e-08, -1.58343e-09, 
    1.463775e-10, 3.996092e-10, -1.018279e-10, 9.351595e-10, -1.235414e-09, 
    1.931198e-09, 2.98968e-09, 1.072506e-08, -7.068195e-10, -1.001695e-09, 
    8.569032e-09, 1.674437e-09, 2.117588e-09, 1.256467e-09, 1.702898e-08, 
    2.689043e-08, 9.003543e-09, -1.129996e-08, 2.852971e-10, -6.355641e-08, 
    4.822368e-09, 3.731161e-08, 1.913456e-10, 2.22276e-08, 7.597123e-10, 
    -5.03178e-11, -2.091667e-09, -3.651017e-10, -6.485919e-09, 1.875893e-09, 
    1.163096e-08, 7.845983e-09, 2.229399e-10, -1.038023e-08, 1.177142e-08, 
    5.768982e-09, -1.036256e-09, -3.863079e-09, 3.786226e-09, -1.942567e-08, 
    -1.641263e-08, -1.61549e-11, 7.859526e-10, -1.478462e-10, -3.69802e-11, 
    -3.112177e-10,
  -8.307666e-10, -9.457608e-10, -1.27875e-09, 6.326673e-11, 3.168736e-09, 
    2.330523e-09, 1.140847e-09, 5.991296e-10, -5.741526e-09, -1.250396e-08, 
    -3.409014e-09, -9.233418e-09, 1.251351e-09, 8.527195e-09, 1.290044e-08, 
    -4.656221e-09, -5.849955e-09, 3.791598e-09, -7.434345e-09, 2.070237e-10, 
    1.707633e-09, 1.612307e-09, 7.435119e-10, 3.176297e-09, -5.473453e-10, 
    1.236344e-10, 6.715254e-08, -1.805472e-08, -1.980635e-08, 2.55244e-09, 
    3.175569e-08, -1.672674e-09, 1.048079e-08, -1.111977e-08, 1.298872e-10, 
    3.877068e-08, -3.34357e-09, 4.125411e-11, -1.506146e-08, -1.527146e-08, 
    -1.28987e-08, 3.914181e-09, -1.36572e-09, -3.308652e-09, -5.297238e-10, 
    -1.235497e-08, -1.539664e-08, -1.933954e-08, -8.74594e-09, -7.301182e-11, 
    -6.327213e-09, -6.602363e-10, 7.962496e-09, 3.797652e-09, 1.328148e-09, 
    1.053877e-10, -4.988817e-08, 1.368477e-09, 3.248327e-08, -1.301196e-08, 
    4.769333e-09, 2.346496e-10, -2.452964e-09, -2.720168e-08, 3.953266e-09, 
    -5.269385e-11, 2.025752e-08, -3.083142e-08, -2.062774e-08, -1.850066e-08, 
    -9.338038e-08, -1.108162e-09, -4.102401e-08, -2.782485e-09, 1.763425e-09, 
    9.693508e-10, -7.667467e-11, 2.092165e-09, -1.576585e-09, 2.008676e-09, 
    3.661143e-09, 1.33183e-08, -6.705534e-10, -3.043397e-10, 1.173589e-09, 
    1.949672e-09, -1.435922e-09, 2.150273e-09, 7.190742e-09, 2.888433e-08, 
    5.216464e-09, -2.09831e-08, -7.998437e-10, -1.053782e-07, 1.194138e-08, 
    -5.898448e-09, 4.06942e-09, 1.704444e-08, -2.30898e-10, -1.277726e-10, 
    -1.626802e-09, -2.386571e-10, -9.168613e-09, 3.092079e-09, 4.185551e-09, 
    1.464514e-09, -6.218272e-09, -7.324275e-10, 9.617906e-09, 1.103501e-09, 
    -5.697416e-10, -4.799858e-09, 4.850619e-09, -6.249195e-09, -1.973177e-08, 
    -1.188027e-12, 8.741665e-10, -1.489582e-10, -4.948575e-11, 7.804601e-11,
  -1.599346e-09, -4.673666e-10, -2.996785e-10, -3.191758e-09, -1.867875e-10, 
    -1.020169e-09, 2.885145e-09, -6.206506e-09, 6.455252e-09, -7.290566e-09, 
    -6.950188e-09, -4.256663e-09, 6.880555e-09, 1.05149e-08, 2.468312e-08, 
    -4.558808e-09, -8.364292e-09, 2.499974e-09, -6.15109e-09, 1.22958e-09, 
    2.053127e-09, 5.887273e-09, -2.13646e-09, 4.321237e-09, -6.70866e-10, 
    8.860752e-10, 7.215749e-08, -3.386765e-08, -2.959939e-08, -5.077595e-09, 
    3.998042e-08, -1.612307e-09, 1.588944e-08, -1.391493e-08, 1.162226e-08, 
    3.512537e-08, -2.192758e-09, 7.915446e-11, -4.073968e-09, -2.092786e-08, 
    -1.1411e-08, 3.104049e-09, -2.547722e-10, -2.752094e-09, 5.171842e-09, 
    2.972439e-08, -1.433838e-08, -2.54048e-08, -1.826891e-08, -1.571863e-10, 
    -4.759912e-09, 2.522484e-09, 1.368101e-08, 5.667641e-09, 1.821951e-09, 
    -6.906475e-12, -5.971253e-08, 1.35272e-09, 3.893027e-08, 3.660716e-11, 
    2.857007e-09, 1.518288e-10, -2.687727e-09, -1.826658e-08, -1.843e-09, 
    3.858418e-09, 2.275465e-08, -2.840892e-08, -3.16918e-08, -1.293824e-08, 
    -1.08983e-07, -3.992966e-09, -5.874955e-08, -3.12383e-09, 4.825307e-09, 
    1.375895e-09, -2.796838e-10, 3.08043e-09, -2.11367e-09, 1.196327e-09, 
    5.957816e-09, 5.349766e-09, -3.269349e-10, 7.889298e-10, -2.321428e-09, 
    2.61025e-10, -5.999766e-09, 5.547236e-09, -5.551721e-09, 2.539085e-08, 
    1.544322e-09, -2.452408e-08, -2.336677e-09, -9.706702e-08, 1.254517e-08, 
    -6.296813e-08, 2.694236e-10, 3.747573e-09, -2.86019e-09, -5.412062e-10, 
    1.523404e-10, -4.414957e-11, -1.34948e-08, 4.814556e-09, 9.757173e-10, 
    -7.956146e-09, -5.846005e-09, 8.069776e-09, 5.786205e-09, 6.118057e-10, 
    3.337846e-10, -2.83751e-09, -2.019078e-09, 7.226902e-09, -6.512948e-09, 
    9.492851e-12, 4.656897e-10, -1.588436e-10, -3.991119e-11, 6.986056e-11,
  -1.470369e-09, -3.791456e-11, 5.246648e-11, -2.633271e-09, -4.015817e-09, 
    -5.135632e-09, -3.249511e-09, -9.762687e-09, 1.862099e-08, 3.009234e-09, 
    1.919432e-09, 3.974264e-09, 3.105413e-09, 5.470213e-09, 2.965277e-08, 
    6.030008e-10, -1.203345e-08, -1.769109e-09, -2.38893e-09, 1.680121e-09, 
    -4.757283e-09, 6.653693e-09, 5.964353e-09, 4.689696e-09, -4.454819e-10, 
    1.096168e-09, -4.86807e-10, -4.291098e-08, -2.71599e-08, -9.184021e-09, 
    4.746659e-08, -7.933124e-09, 2.484063e-08, -3.085972e-09, 1.228892e-08, 
    3.008427e-08, -9.259736e-10, 1.619327e-10, 4.779224e-09, -2.784201e-08, 
    -3.619266e-09, -2.577281e-10, 3.101889e-09, 1.980237e-08, 4.525566e-08, 
    4.99117e-08, -1.373212e-08, -3.206466e-08, -2.62021e-08, -2.463274e-10, 
    -5.702411e-09, 3.36513e-09, 2.221731e-08, 8.664472e-09, 2.845222e-09, 
    -1.147384e-10, -6.033594e-08, 2.964134e-09, -1.474285e-08, 1.122935e-09, 
    -3.779348e-09, -2.530726e-09, -3.402874e-09, -4.481035e-09, 
    -8.521374e-09, 6.796711e-09, 2.210385e-08, -1.800436e-08, -4.132067e-08, 
    -7.725362e-09, -9.048478e-08, -2.246281e-09, -7.409761e-08, 
    -3.013497e-09, 3.860896e-09, 1.859576e-09, -2.279066e-10, 3.214112e-09, 
    -2.337105e-09, 9.068799e-10, 1.075585e-08, -6.896052e-09, 3.383889e-10, 
    1.314163e-09, -1.711953e-09, -2.169827e-09, -7.943868e-09, 7.18029e-09, 
    -1.804016e-08, 1.610096e-08, -3.640821e-10, -2.716309e-08, -3.31049e-09, 
    -7.806786e-08, 2.021892e-08, -7.040401e-08, 6.141988e-09, 9.295206e-09, 
    -5.656204e-09, -1.744149e-09, 1.875037e-09, 5.199112e-10, -2.096798e-08, 
    7.677972e-09, -1.177341e-09, -6.764992e-09, 4.980166e-09, 1.059357e-08, 
    2.806303e-09, 6.615437e-10, 2.444267e-10, -3.832952e-10, -2.956256e-09, 
    9.425491e-09, 1.06017e-08, 2.914362e-11, 7.312195e-11, -1.431371e-10, 
    5.610801e-11, -1.979288e-10,
  -2.512479e-10, 1.98952e-11, 3.32841e-09, 4.478352e-09, -6.148412e-09, 
    -4.175376e-09, -9.341875e-09, -8.690904e-09, 1.508693e-08, 1.650346e-08, 
    1.310673e-08, 5.612719e-09, 2.039542e-10, 1.051717e-09, 8.270376e-09, 
    1.266202e-08, -2.001041e-08, -5.518018e-09, 1.422976e-09, 1.673243e-09, 
    -2.758202e-08, -4.195613e-08, -3.107482e-08, -3.880359e-09, 5.892389e-10, 
    8.385541e-10, 3.103651e-11, -4.120113e-08, -4.2946e-08, -1.685032e-08, 
    4.036099e-08, -1.446119e-08, 3.446019e-08, 4.906724e-10, 7.76879e-09, 
    4.545018e-08, -1.321223e-09, 1.865885e-10, 2.201796e-08, -3.620763e-08, 
    1.147464e-09, -8.416237e-10, 5.181619e-09, 2.249791e-08, 4.061633e-08, 
    1.855574e-08, -1.357284e-08, -4.47935e-08, -3.104033e-08, -2.593907e-10, 
    -3.42817e-09, 1.078172e-08, 2.086079e-08, 9.996734e-09, 4.206854e-09, 
    -3.138325e-10, -4.949618e-08, 9.982795e-09, -4.437519e-08, -6.332073e-10, 
    -9.594032e-10, -4.79497e-09, -1.336389e-09, 1.242975e-08, -1.404551e-08, 
    6.328264e-09, 1.247645e-08, -2.570573e-09, -1.981812e-08, -7.308472e-09, 
    -9.350822e-08, -1.329579e-08, -5.838399e-08, 1.789999e-09, -3.858338e-09, 
    2.787147e-09, 3.261533e-10, 2.286953e-09, -2.062626e-09, 4.218919e-10, 
    1.824014e-08, -4.191457e-09, 9.541736e-10, 4.498588e-10, -2.694037e-09, 
    1.042281e-09, -1.319063e-08, 6.145342e-09, -2.657691e-08, -7.244694e-10, 
    -2.232696e-09, -2.570857e-08, -3.720345e-09, -1.235833e-08, 1.748936e-08, 
    -1.378894e-08, 1.151968e-08, 2.789886e-08, -7.72593e-09, -3.805281e-09, 
    1.554213e-09, -1.320345e-09, -2.938148e-08, 9.768584e-09, -4.70834e-09, 
    -6.259711e-09, -4.962089e-09, 5.401489e-09, 9.403038e-10, -7.833023e-10, 
    -1.370267e-09, -4.539515e-10, -1.740887e-09, 7.286417e-09, 1.488252e-08, 
    1.442686e-11, -6.542678e-11, -1.440519e-10, 9.475087e-11, 5.625225e-10,
  -9.396217e-11, 5.553602e-11, 5.12847e-09, 2.285589e-08, -3.170669e-09, 
    -3.208982e-09, -8.901054e-09, -3.357115e-09, -1.737646e-09, 1.783013e-08, 
    1.403799e-08, 1.164722e-10, -1.520277e-09, -7.48571e-10, -7.054837e-10, 
    3.20394e-08, -2.988571e-08, -3.201876e-09, 4.369184e-09, -2.924423e-09, 
    -5.665089e-08, -5.970566e-08, -5.906981e-08, -1.061886e-08, 1.632372e-09, 
    1.221395e-09, -1.503525e-08, -2.565929e-08, -5.040766e-08, -1.952395e-08, 
    2.03915e-08, -3.391102e-08, 4.543978e-08, 9.477333e-09, 2.476611e-09, 
    4.325494e-08, -1.959188e-09, 1.706724e-10, 1.446057e-08, -4.055016e-08, 
    -9.683507e-10, 1.739124e-09, 3.535661e-09, 1.421328e-08, 8.642417e-09, 
    1.624443e-08, -1.257553e-08, -5.780629e-08, -3.586593e-08, -3.324914e-10, 
    1.930175e-09, 9.746657e-09, 1.010101e-08, 1.145785e-08, 4.258453e-09, 
    -4.801564e-10, -3.256304e-08, 1.754753e-08, -2.023801e-08, -8.690193e-09, 
    7.254869e-09, -2.44296e-09, 2.158345e-10, 8.851191e-09, -2.299982e-08, 
    1.200073e-08, -2.927436e-11, 1.535312e-08, 1.796792e-08, -4.870742e-09, 
    -1.240711e-07, -3.202314e-08, -5.911016e-08, 4.580841e-09, -3.362908e-08, 
    2.035165e-09, -9.583374e-10, 1.384024e-09, -2.124725e-09, 1.066951e-10, 
    2.359405e-08, 3.524875e-08, 1.146134e-09, -2.56199e-09, -6.98094e-10, 
    7.322171e-09, 1.300634e-09, 3.624734e-09, -2.746209e-08, -1.844967e-08, 
    -4.360743e-09, -2.207552e-08, -3.528982e-09, 5.720159e-08, 5.926665e-09, 
    1.626377e-08, 1.196464e-08, 2.05377e-08, -9.758594e-09, -6.01766e-09, 
    -1.281649e-09, -1.54048e-08, -2.483824e-08, 8.929284e-09, -3.039474e-09, 
    -9.856137e-09, -1.792199e-08, 1.044197e-08, 2.721379e-09, -1.91659e-09, 
    -2.246281e-09, -1.351168e-10, 1.214744e-10, 2.247873e-09, 4.208744e-09, 
    1.529088e-10, -2.99238e-10, -5.851319e-11, 1.824958e-10, 3.873708e-09,
  4.495519e-09, 2.972911e-10, 2.415618e-09, 2.471279e-08, 6.993218e-09, 
    -1.648459e-11, -7.703647e-09, -8.960797e-10, -1.393755e-08, 6.035521e-09, 
    7.818926e-09, -1.905619e-09, -2.377192e-09, -1.662136e-08, -1.985768e-09, 
    5.140363e-08, -4.108107e-08, -4.258538e-09, 8.310749e-09, -1.184628e-08, 
    -6.528614e-08, -3.62927e-08, -3.431671e-08, -1.926571e-08, 1.478043e-09, 
    1.815238e-09, -9.887003e-09, -2.245702e-08, -2.872059e-08, 2.939373e-09, 
    -2.274589e-08, -4.651099e-08, 5.473782e-08, -2.896059e-09, -4.71664e-09, 
    1.791e-08, -7.071662e-10, 4.126832e-11, -1.285628e-08, -3.958191e-08, 
    -7.119934e-09, 2.359002e-09, 5.672973e-10, 5.967793e-09, 9.964651e-09, 
    -9.966925e-10, -1.039677e-08, -6.846417e-08, -3.151863e-08, 
    -2.148248e-09, 1.298103e-08, 4.336925e-09, 7.454332e-09, 1.417734e-08, 
    1.999666e-09, -5.022684e-10, -1.11437e-08, 3.150836e-08, 1.066819e-08, 
    -1.092968e-08, 8.712959e-09, -2.349907e-10, 1.467697e-10, 4.523144e-10, 
    -3.678824e-08, 3.06876e-08, -8.014354e-09, 2.514694e-07, 3.082266e-08, 
    5.85635e-09, -1.827631e-07, -4.07789e-08, -4.478488e-08, 2.551019e-09, 
    -7.288546e-08, -1.241233e-09, -1.055682e-09, -9.646328e-11, 
    -1.788433e-09, -5.705942e-10, 2.488076e-08, 9.432569e-08, 8.660663e-10, 
    -4.841468e-09, 1.270337e-09, 1.147657e-08, 2.123272e-08, 1.658805e-09, 
    -2.113593e-08, -3.291319e-08, -4.966523e-09, -2.186132e-08, 
    -1.963059e-09, 1.104396e-07, 1.046317e-08, 5.52069e-08, 1.637297e-09, 
    2.054912e-08, -1.055525e-08, -7.720178e-09, -1.570993e-08, -3.422166e-08, 
    -1.733005e-08, 5.3479e-09, -3.069886e-09, -1.60386e-08, -2.354432e-08, 
    1.940998e-08, 8.845177e-09, -5.528591e-10, -2.226784e-09, 1.297849e-09, 
    4.844196e-10, -6.3568e-09, -2.442562e-09, 6.112146e-10, -2.735447e-10, 
    2.04281e-11, 2.880185e-10, 7.807216e-09,
  3.499963e-08, 1.695071e-10, 4.370122e-10, 9.770815e-09, 1.635351e-08, 
    1.035164e-08, -7.901008e-09, -2.616162e-09, -3.758032e-09, -1.090064e-08, 
    -4.219032e-09, -5.033598e-09, -1.455192e-11, -5.159541e-08, 4.649792e-11, 
    7.022777e-08, -5.265318e-08, -9.753649e-09, 2.098764e-08, -2.299191e-08, 
    -3.337266e-08, -2.24702e-08, -6.414211e-10, -1.193973e-08, 3.061814e-09, 
    8.358256e-10, 2.757973e-07, -2.874162e-08, -5.877723e-09, 7.685969e-08, 
    3.527362e-09, -3.149512e-08, 6.937228e-08, 7.106678e-09, -3.536331e-08, 
    -1.145679e-08, 3.424725e-09, -2.07649e-10, -4.630954e-08, -4.626236e-08, 
    -1.896908e-08, 8.880079e-10, -3.566072e-10, -6.305195e-09, 4.170693e-08, 
    -1.493868e-08, -7.533288e-09, -8.356477e-08, -2.29981e-08, 4.607017e-10, 
    2.228768e-08, -1.487717e-08, 1.626175e-08, 1.836465e-08, -4.219231e-10, 
    -5.667289e-11, 5.846459e-09, 5.379013e-08, 7.237225e-09, -1.444702e-08, 
    3.721084e-09, 2.728484e-11, 1.210765e-10, 1.617127e-09, -5.353197e-08, 
    9.065434e-08, -1.884143e-08, 2.002198e-07, 3.08612e-08, -1.861952e-08, 
    -2.420988e-07, -3.45027e-08, -2.608738e-08, 2.554657e-09, -7.834316e-08, 
    -9.082328e-09, 1.83519e-10, -3.390312e-09, -1.53596e-09, -2.577622e-09, 
    1.339237e-08, 1.170376e-07, 1.357989e-10, -5.371476e-09, -7.752305e-09, 
    1.167018e-08, 2.051183e-08, 5.045422e-10, -1.14206e-08, -3.074308e-08, 
    -1.920284e-09, -1.687006e-08, 7.782432e-10, 1.715444e-07, 8.867573e-09, 
    9.096004e-08, -1.155238e-08, 2.315426e-08, -1.575131e-08, -9.409336e-09, 
    -3.441846e-08, -4.433371e-08, -1.104738e-08, 3.391065e-09, 5.794277e-09, 
    -1.922206e-08, -2.972945e-08, 3.298805e-08, 1.639785e-08, 8.143388e-10, 
    -3.898322e-10, 2.410388e-09, -2.989623e-09, -1.502337e-08, -3.722107e-10, 
    9.530594e-10, 3.009859e-11, -7.979395e-12, 3.657235e-10, 1.534431e-08,
  6.604137e-08, 1.477929e-11, 1.121066e-09, 1.041394e-08, 3.520336e-08, 
    2.427464e-08, -5.049174e-09, -4.569984e-09, -3.004402e-09, -3.397076e-09, 
    -8.624397e-09, -1.104195e-08, -5.960601e-10, -6.554785e-08, 2.497131e-09, 
    8.492778e-08, -6.567321e-08, -1.148771e-08, 3.766496e-08, -4.189587e-08, 
    1.888191e-08, -2.885645e-08, 1.075364e-08, -3.608989e-09, -5.437641e-10, 
    -8.092229e-10, 3.486437e-07, -2.409035e-08, -1.042247e-08, 1.461821e-07, 
    -1.988531e-08, -3.892148e-08, 6.61779e-08, 2.317273e-07, -6.835364e-08, 
    -8.06773e-08, 5.922402e-10, -6.852332e-10, -6.074004e-08, -4.409488e-08, 
    -3.71125e-08, 7.914878e-10, -3.500875e-08, -1.466542e-08, 6.922517e-08, 
    1.627836e-08, -6.608843e-09, -1.012079e-07, -1.904123e-08, 1.008198e-08, 
    3.269416e-08, -2.522427e-08, 3.485599e-08, 2.424531e-08, -4.615759e-09, 
    -2.638103e-10, 1.983528e-08, 9.519296e-08, -9.185535e-08, -1.595009e-08, 
    1.706212e-09, -4.562253e-10, -2.064553e-10, 2.361662e-08, -6.703299e-08, 
    7.707945e-08, -5.693141e-08, 5.439301e-08, -4.447088e-09, -9.007863e-09, 
    -2.39648e-07, -4.301114e-08, -1.577826e-08, 1.228227e-08, -3.471198e-08, 
    -2.484512e-09, 2.811191e-10, -5.170961e-09, -1.086201e-09, -1.279045e-07, 
    -5.417178e-09, 9.852439e-08, -8.654979e-10, -6.725941e-09, -1.551928e-08, 
    -2.686318e-08, -3.80976e-09, 1.192234e-09, -7.428227e-09, -1.991299e-08, 
    1.790568e-09, -8.676693e-09, 3.039304e-09, 2.308747e-07, 2.375032e-09, 
    1.031229e-07, -1.426863e-08, 1.641323e-07, -2.438685e-08, -1.136161e-08, 
    -1.221258e-08, -4.412082e-08, -5.774012e-09, 1.790035e-09, -1.429623e-08, 
    -2.05182e-09, -9.202722e-09, 3.17026e-08, 2.519459e-08, 6.386927e-10, 
    3.145374e-09, 8.005827e-10, -7.442395e-09, -1.303249e-08, 1.754188e-10, 
    7.239237e-10, 3.425384e-10, 9.718804e-11, 4.05727e-10, 1.924263e-08,
  5.82163e-08, -1.20508e-11, 2.631396e-09, 2.420836e-08, 3.710863e-08, 
    2.982881e-08, -1.118678e-10, -6.27233e-09, -1.316141e-08, -1.140154e-08, 
    -4.838398e-09, -6.374648e-09, -3.148784e-09, -4.639571e-08, 3.197215e-09, 
    8.755279e-08, -8.02158e-08, -1.474422e-08, 5.641202e-08, -7.595906e-08, 
    6.276514e-08, -5.513914e-08, 8.819825e-10, -3.284526e-09, -9.338237e-09, 
    4.24734e-10, 7.753101e-09, -1.545266e-08, -4.160825e-09, 6.212383e-08, 
    -7.514132e-09, -4.997435e-08, 5.085656e-08, 3.216894e-07, -8.456766e-08, 
    -1.187228e-07, -9.304699e-09, -9.544436e-10, -5.457366e-08, 
    -3.611049e-08, -4.836081e-08, 2.707338e-09, -1.472874e-07, -2.340466e-08, 
    3.475304e-08, 5.290656e-08, -1.545953e-08, -1.199701e-07, -1.526191e-08, 
    2.073466e-08, 3.943498e-08, -7.656149e-08, 5.704133e-08, 2.869663e-08, 
    -7.664485e-09, -8.299708e-10, 3.36006e-08, 1.379685e-07, -1.76926e-07, 
    -1.940644e-08, 3.558512e-09, -4.214371e-10, 6.286882e-11, 4.604354e-08, 
    -7.537437e-08, 1.365418e-07, -9.141229e-08, -2.039974e-08, -6.654318e-09, 
    -3.816467e-10, -2.614097e-07, -5.335346e-08, -1.118576e-08, 2.014781e-08, 
    -2.756769e-09, -2.053525e-09, 5.078959e-11, -4.080817e-09, -8.993226e-10, 
    -2.283314e-07, -1.726858e-08, 5.926941e-08, -1.349292e-09, 1.724402e-09, 
    -9.560608e-09, -8.653387e-08, 2.797361e-07, 1.738158e-09, -1.081366e-08, 
    -9.019573e-09, 2.974048e-09, 3.076366e-10, 3.8861e-09, 2.326068e-07, 
    -1.588296e-08, 1.200066e-07, 5.108497e-09, 7.313645e-08, -4.191975e-08, 
    -1.249509e-08, 4.859555e-08, -2.754737e-08, -7.44469e-09, 1.422698e-09, 
    -6.930577e-08, 2.27293e-08, 2.55227e-10, 3.075138e-08, 3.545745e-08, 
    -3.237801e-10, 2.986894e-09, -1.365379e-10, -9.513656e-09, -9.454993e-09, 
    -1.759076e-09, 8.982397e-10, -1.008971e-12, -2.9587e-10, 4.406289e-10, 
    1.412411e-08,
  3.402209e-08, 2.12026e-11, 8.266227e-09, 3.421286e-08, 3.263136e-08, 
    2.591133e-08, 1.048136e-09, -4.815945e-09, -1.439838e-08, -1.607702e-09, 
    -3.332673e-09, 5.974243e-11, -9.524626e-09, 4.662809e-09, 5.083564e-09, 
    7.678477e-08, -8.808333e-08, -2.344615e-08, 7.805654e-08, -1.289944e-07, 
    8.256876e-08, -6.758438e-08, -3.127468e-09, -3.515254e-09, -3.913044e-09, 
    5.020468e-09, -2.267626e-08, -9.782582e-09, -2.330182e-09, -1.717564e-08, 
    2.743661e-09, -2.856456e-08, 2.894586e-08, 1.673885e-07, -7.876423e-08, 
    -6.109548e-08, -2.053152e-08, -1.185029e-09, -6.03381e-08, -2.264023e-08, 
    -4.574318e-08, 2.467289e-09, -1.284556e-07, -3.446843e-08, 1.810344e-08, 
    6.750275e-08, -1.676761e-08, -1.38351e-07, -9.881058e-09, 2.711622e-08, 
    4.34964e-08, -1.414695e-07, 6.258199e-08, 3.433957e-08, -1.124196e-08, 
    -1.474916e-09, 4.475015e-08, 1.759289e-07, -2.874101e-07, -2.857595e-08, 
    4.610968e-09, 1.956948e-09, -2.086153e-11, 6.383819e-08, -8.236749e-08, 
    1.447268e-07, -7.898615e-08, 8.510489e-08, 2.249641e-08, 9.670487e-09, 
    -2.718935e-07, -3.396195e-08, -2.55389e-08, 1.477264e-08, 1.063204e-08, 
    -1.9531e-08, -9.40247e-10, 1.337099e-09, -4.327455e-09, -1.602444e-07, 
    -2.466629e-08, 1.826427e-08, 4.039862e-10, 9.117286e-09, 8.283791e-10, 
    -2.934547e-08, 2.065082e-08, 1.974342e-09, -2.334097e-08, 5.38023e-10, 
    1.934382e-10, 2.963601e-09, 5.500738e-09, 2.054399e-07, -1.827738e-08, 
    1.443116e-07, 4.944321e-08, 1.597215e-08, -5.812302e-08, -1.140298e-08, 
    7.30509e-08, 2.257899e-09, -1.302209e-08, 7.929515e-10, -8.25541e-08, 
    -7.164829e-09, -6.443486e-09, 2.544931e-08, 5.805515e-08, -2.686988e-10, 
    1.202523e-09, 4.818901e-09, -9.562143e-09, -5.906202e-09, 7.333369e-10, 
    1.594287e-09, -1.06462e-09, -9.140315e-10, 5.254464e-10, -1.729853e-08,
  1.508602e-08, -5.84123e-10, 9.377118e-09, 2.637807e-08, 2.271952e-08, 
    1.655349e-08, -6.199343e-10, -2.364686e-09, -8.163738e-09, 8.137704e-10, 
    6.780738e-09, 1.607418e-09, -7.825633e-09, 1.179137e-08, 1.865499e-08, 
    5.11342e-08, -8.007174e-08, -2.989128e-08, 1.011592e-07, -1.464201e-07, 
    5.853633e-08, -5.009178e-08, -4.291905e-09, -1.788976e-09, 4.253366e-09, 
    4.730782e-08, -3.315552e-08, -1.049466e-08, 5.243919e-09, -4.750291e-09, 
    3.435389e-09, -1.058254e-08, 2.142087e-08, -1.408757e-07, -7.155268e-08, 
    -1.443675e-08, -3.7733e-08, -2.379494e-09, -8.705069e-08, -4.087376e-09, 
    -2.792376e-08, 9.066525e-10, -1.715327e-08, -2.923844e-08, 2.110755e-08, 
    8.092627e-08, -1.385609e-08, -1.556058e-07, -1.020214e-08, 3.080844e-08, 
    4.39685e-08, -1.65626e-07, 4.478927e-08, 3.802727e-08, -1.490023e-08, 
    8.084839e-10, 5.393042e-08, 1.131409e-08, -3.731579e-07, -5.192223e-08, 
    3.258151e-09, 2.887293e-08, -4.429614e-08, 7.789109e-08, -9.130345e-08, 
    3.952596e-08, -7.724964e-08, 8.918437e-08, 2.468528e-08, 2.260322e-08, 
    -1.719676e-07, -1.495391e-08, -4.504409e-08, 2.914589e-09, 1.271314e-08, 
    -2.280694e-08, 1.284448e-09, 9.572062e-09, -4.721528e-09, -5.489142e-08, 
    -3.680373e-08, -2.991035e-09, 4.445326e-09, 6.189566e-09, -2.109914e-09, 
    -4.413891e-09, -1.692949e-07, -6.161827e-11, -3.148503e-08, 2.240029e-09, 
    8.726829e-09, 1.524176e-09, 7.217238e-09, 1.762989e-07, -9.353926e-09, 
    1.800674e-07, 9.31487e-08, 3.391892e-08, -7.175288e-08, -9.097743e-09, 
    -7.558697e-09, 2.284471e-08, -5.517698e-09, 8.169678e-10, -9.91605e-08, 
    -2.83851e-08, 2.018169e-08, -4.270646e-09, 7.79653e-08, -9.030146e-10, 
    6.286882e-11, 1.524643e-08, -2.361389e-09, -4.17117e-10, 3.728246e-09, 
    2.304114e-09, -3.198522e-09, -9.847341e-10, 6.114718e-10, -3.522439e-08,
  7.281756e-09, -6.272899e-09, 7.983431e-09, 3.478476e-09, 1.104706e-08, 
    1.041565e-08, -3.081482e-09, 6.494588e-09, -8.022766e-09, -5.254049e-08, 
    8.177494e-10, 1.169269e-09, -5.330833e-08, -4.675337e-08, 4.549713e-08, 
    1.193571e-08, -5.968013e-08, -3.564423e-08, 1.176416e-07, -8.963173e-08, 
    1.085971e-08, -1.849378e-08, -7.511403e-09, -8.695906e-10, -1.214744e-09, 
    1.21105e-07, -3.064622e-08, 1.572073e-08, 1.337264e-08, 8.838128e-09, 
    1.058027e-08, -1.245439e-09, 2.887248e-08, -8.124482e-08, -6.653488e-08, 
    1.182286e-08, -5.552938e-08, -2.478885e-09, -1.266313e-07, 1.659682e-08, 
    1.312226e-08, -1.614012e-09, 7.277237e-08, -2.1468e-08, 1.368846e-08, 
    6.854305e-08, -6.155346e-09, -1.710139e-07, -1.015576e-08, 2.972192e-08, 
    4.165037e-08, -1.873381e-07, 2.462511e-08, 4.794613e-08, -1.766217e-08, 
    4.835101e-10, 5.835989e-08, 1.482404e-07, -3.975286e-07, -5.797861e-08, 
    2.179945e-09, 5.891263e-08, -1.3072e-07, 1.174918e-07, -9.797448e-08, 
    6.364701e-08, -6.454241e-08, -4.233129e-09, 3.246328e-09, 2.812578e-08, 
    -3.174171e-08, -3.631726e-09, -4.076321e-08, -2.662432e-09, 4.70518e-09, 
    -1.911383e-08, 3.483478e-09, 2.042083e-08, -7.560686e-10, -4.524384e-08, 
    -6.91681e-08, -3.333622e-09, 9.967835e-09, -3.807656e-08, 2.216552e-09, 
    -1.304045e-08, -9.077792e-08, -3.863875e-09, -4.255884e-08, 
    -8.952952e-09, 1.997535e-08, -4.268781e-09, 4.491937e-09, 2.063377e-07, 
    -9.921337e-09, 1.848332e-07, 1.521697e-07, 1.881983e-08, -8.562586e-08, 
    -9.763949e-09, -3.752803e-10, 1.25589e-08, -1.032953e-08, 5.554597e-10, 
    -8.702762e-08, 2.930381e-08, 3.544017e-08, -1.149635e-08, 7.43006e-08, 
    -3.326363e-09, -1.817284e-09, 2.154695e-08, 1.632372e-08, 1.608669e-10, 
    1.015565e-09, 2.907996e-09, -1.81339e-09, -1.014278e-09, 6.511414e-10, 
    -1.337742e-08,
  6.826156e-09, -2.282633e-08, 2.617924e-09, -3.4572e-08, -5.917002e-09, 
    4.320498e-09, 1.94575e-10, 1.757456e-08, -6.918583e-09, -9.858405e-08, 
    -4.258692e-08, -1.863629e-08, -5.670091e-08, -1.05589e-07, 2.081282e-08, 
    -1.067281e-09, -3.167776e-08, -4.271539e-08, 1.221792e-07, -7.510891e-09, 
    -8.178233e-09, 9.503253e-09, -1.184168e-08, -2.369802e-10, 1.062034e-08, 
    1.448965e-07, -2.520466e-08, 2.403129e-08, 1.775646e-08, 4.802968e-08, 
    1.164371e-07, -4.086473e-10, 4.308384e-08, -2.972894e-08, -4.185205e-08, 
    3.19987e-08, -6.079264e-08, -2.672778e-09, -1.400804e-07, 3.016864e-08, 
    3.940903e-08, -1.70615e-08, 2.416436e-08, -1.389364e-08, 8.482118e-09, 
    4.181646e-08, 2.276812e-08, -1.83762e-07, -1.162535e-08, 2.324926e-08, 
    3.832358e-08, -2.182554e-07, 1.293435e-08, 6.01908e-08, -2.20703e-08, 
    9.261498e-10, 6.242698e-08, 2.242029e-07, -4.870736e-07, -3.757239e-08, 
    2.107697e-09, -3.669976e-08, -1.890906e-07, 1.600001e-07, -1.004629e-07, 
    6.21128e-10, -4.195527e-08, -3.671499e-08, 1.769666e-08, 2.271207e-08, 
    5.570558e-08, 2.016867e-08, -2.644157e-08, -6.06093e-09, 3.702132e-09, 
    -1.798441e-08, 8.7648e-09, 3.408002e-08, -2.669765e-09, -1.039883e-07, 
    -1.10608e-07, -5.14301e-09, 1.038194e-08, -9.205434e-08, -2.183384e-08, 
    -1.881136e-08, -9.790284e-08, -1.271587e-10, -7.103058e-08, 
    -2.958399e-08, 3.257526e-09, -1.030813e-08, 2.818979e-09, 2.275102e-07, 
    1.101597e-08, 1.945979e-07, 1.863752e-07, -7.033242e-08, -9.46464e-08, 
    -9.913685e-09, 8.904578e-09, -1.499333e-08, -1.876273e-08, 4.864944e-09, 
    -8.208195e-08, 9.080048e-08, -4.528766e-08, -5.584127e-09, 4.25627e-08, 
    -6.725543e-09, -1.117911e-08, 1.640495e-08, 3.240433e-08, 9.144401e-10, 
    -1.068412e-08, 3.386833e-09, -2.551786e-09, -8.730723e-10, 7.847092e-10, 
    -2.938378e-08,
  1.060727e-08, -4.624229e-08, 1.874298e-09, -5.032547e-08, -4.466159e-08, 
    -6.979803e-10, 5.022741e-09, 2.233543e-08, -8.409984e-10, -6.622457e-08, 
    -6.267277e-08, -2.422297e-08, -1.709981e-08, -7.751549e-08, 8.304823e-11, 
    4.159131e-09, -2.886804e-08, -3.237943e-08, 8.693524e-08, 1.698143e-07, 
    -3.854067e-07, 3.316529e-09, -5.880963e-09, 1.420688e-09, 3.934434e-08, 
    9.201318e-08, -4.712717e-09, 2.465623e-08, 1.410245e-08, 1.94637e-08, 
    1.690117e-07, -2.370433e-08, 1.941413e-08, -1.345231e-07, -2.649534e-08, 
    8.131002e-08, -4.889749e-08, -4.03395e-09, -1.401192e-07, 3.264412e-08, 
    3.211672e-08, -2.546739e-08, -8.642627e-08, -1.027492e-08, 1.30363e-08, 
    2.584153e-08, 2.352905e-07, -1.758559e-07, -2.408755e-08, 1.395011e-08, 
    3.575565e-08, -2.587412e-07, -4.773062e-09, 6.82494e-08, -2.84246e-08, 
    1.012552e-09, 7.704926e-08, 1.991323e-07, -6.237469e-07, -2.620618e-08, 
    5.525749e-10, -6.29372e-08, -1.59265e-07, 1.652998e-07, -8.709802e-08, 
    3.726865e-08, -4.325324e-08, -3.991153e-08, -7.167444e-09, 3.423776e-08, 
    1.026991e-07, 4.022678e-08, 2.130578e-07, -8.22223e-09, 2.898027e-09, 
    -1.608913e-08, -5.811017e-09, 3.888414e-08, -7.099697e-09, -1.665011e-07, 
    -1.532241e-07, -3.167685e-09, 9.379789e-09, 5.859704e-09, -5.195869e-08, 
    2.589223e-08, -5.306828e-08, 9.146618e-09, -8.860457e-08, -5.316446e-08, 
    1.791869e-08, -1.255197e-08, -6.096798e-09, 2.536183e-07, 1.955556e-08, 
    2.22271e-07, 1.605789e-07, -4.859197e-08, -1.171579e-07, -6.800189e-09, 
    1.564518e-08, -7.082218e-08, -2.46928e-08, 9.824944e-09, -1.108701e-07, 
    4.944337e-08, -1.023481e-07, 5.273364e-10, -3.36621e-09, -1.355937e-08, 
    -3.191866e-08, 5.852883e-09, 2.296093e-08, 2.538201e-08, -1.54734e-08, 
    2.821537e-09, -1.840021e-09, -5.514025e-10, 9.574705e-10, -4.834664e-08,
  1.766551e-08, -6.11347e-08, 8.862969e-09, 1.419551e-09, -4.672489e-08, 
    -2.351101e-09, 1.039854e-08, 1.78332e-08, 1.051109e-08, -2.912105e-08, 
    -5.258147e-08, 8.971767e-09, -1.979396e-08, -3.28709e-08, -9.88581e-09, 
    1.22516e-08, -3.404963e-08, -1.625892e-09, 9.534823e-08, 8.395278e-08, 
    -3.471969e-07, -4.055556e-08, 6.874055e-07, 1.365268e-07, 4.702332e-08, 
    8.391447e-08, 1.116024e-08, 2.490248e-08, 8.854215e-09, 1.318256e-09, 
    5.97642e-08, -7.922978e-08, 5.363171e-08, -8.29811e-08, -2.608755e-08, 
    2.279318e-07, -2.372118e-08, -4.564896e-09, -1.270216e-07, 1.671246e-08, 
    -1.432899e-08, -4.048462e-08, -1.49759e-07, -8.400738e-09, -1.309689e-08, 
    1.11267e-08, 2.562644e-07, -1.582239e-07, -1.172197e-08, 5.342493e-09, 
    3.477702e-08, -2.529069e-07, -1.82379e-08, 7.054283e-08, -3.597721e-08, 
    7.636345e-10, 9.687773e-08, 1.682623e-07, -6.760777e-07, -2.341388e-08, 
    -1.450701e-09, 2.009039e-07, -8.702017e-08, 1.29962e-07, -4.003408e-08, 
    5.622945e-08, -5.116857e-08, -1.536608e-08, -1.011534e-08, 3.885117e-08, 
    9.346417e-08, 2.885457e-08, 1.209136e-07, -1.744985e-08, -7.701217e-09, 
    -4.965216e-09, -1.141784e-08, 4.062619e-08, -1.259758e-08, -2.523007e-07, 
    -1.949348e-07, -1.755302e-09, -1.993158e-09, 1.00751e-08, -7.85347e-08, 
    1.26791e-08, -2.807766e-07, 1.909979e-08, -9.081535e-08, -9.492237e-08, 
    4.869236e-08, -9.039889e-09, -1.748748e-08, 2.820952e-07, 1.204222e-08, 
    2.318397e-07, 1.370828e-07, -5.000476e-08, -1.344254e-07, 2.737477e-09, 
    1.557038e-08, -1.078401e-07, -3.33147e-08, 9.207554e-09, -2.733458e-08, 
    1.394204e-08, -8.022351e-08, 9.638939e-10, -3.236636e-08, -2.742667e-08, 
    -4.845793e-08, 2.888214e-10, 6.247717e-09, 5.535088e-08, -8.851941e-09, 
    6.889536e-10, 3.701075e-10, -6.266205e-10, 1.078398e-09, 2.075541e-08,
  1.355289e-08, -5.228634e-08, 8.258041e-09, 6.705778e-08, 1.065206e-08, 
    2.276295e-09, 1.221684e-08, 1.407108e-08, 2.98449e-08, -1.922388e-09, 
    -2.850487e-08, 3.219225e-07, -2.278597e-08, -2.71279e-08, -1.738971e-08, 
    2.331207e-08, -3.988742e-08, 2.166126e-08, 4.185929e-08, -4.087445e-08, 
    3.54533e-08, 4.960822e-08, 1.64876e-08, 1.916813e-07, 1.033896e-07, 
    1.797594e-07, 2.041639e-08, 2.207167e-08, -3.629054e-09, 7.272257e-08, 
    -2.275323e-08, -3.316194e-08, 1.079532e-07, -2.856666e-09, -1.598249e-08, 
    1.376528e-07, -4.018591e-09, -5.459441e-09, -1.170801e-07, -1.415486e-08, 
    -2.818477e-08, 3.982628e-07, -1.593856e-07, -7.034572e-09, -1.010693e-08, 
    1.090876e-08, 1.061254e-07, -1.107633e-07, -2.125902e-08, -2.177529e-10, 
    3.540518e-08, -1.393613e-08, -2.26832e-08, 7.826844e-08, -4.371999e-08, 
    4.600338e-10, 1.064735e-07, 1.459353e-07, -6.52717e-07, 8.860553e-09, 
    -7.680114e-10, 3.039787e-08, -3.75623e-08, 7.308287e-08, 5.004871e-09, 
    5.581552e-08, -5.08557e-08, 5.32674e-09, 3.886328e-09, 4.300233e-08, 
    8.554372e-08, 3.710517e-08, 1.360587e-08, -4.579982e-08, 1.330987e-08, 
    4.676679e-09, -8.922996e-09, 2.582726e-08, -1.351022e-08, -2.531883e-07, 
    -2.344314e-07, 8.927577e-09, -4.260988e-08, -8.736777e-09, -8.784303e-08, 
    -3.973781e-08, -1.485309e-07, 2.702751e-08, -8.207178e-08, -1.245642e-07, 
    1.123372e-07, -2.426458e-08, -1.444437e-08, 2.693859e-07, 5.053022e-08, 
    2.522846e-07, 1.06915e-07, -7.021339e-08, -1.336177e-07, 2.618765e-09, 
    1.83382e-08, -1.080436e-07, -4.048584e-08, 1.708102e-09, -2.96647e-08, 
    -1.126449e-08, -2.734822e-08, 3.784692e-09, -4.353745e-08, -4.092016e-08, 
    -3.62474e-08, -3.893518e-08, 1.446153e-09, 7.044542e-08, -3.921684e-09, 
    -1.269916e-09, 1.97798e-09, -8.009096e-10, 1.09614e-09, 1.45011e-07,
  5.194579e-09, -2.758225e-08, -8.530151e-09, 8.194434e-08, 7.638005e-08, 
    8.3553e-09, 4.098638e-09, 2.570141e-08, 3.373998e-08, 2.000638e-08, 
    1.371222e-08, 5.030915e-07, -1.78361e-08, -5.114202e-08, 2.103025e-08, 
    2.46479e-08, -1.047812e-08, 6.998982e-08, 7.861701e-09, -1.932476e-07, 
    -1.738044e-09, 1.782275e-07, -1.415708e-07, 5.921265e-08, 1.145938e-07, 
    1.695159e-07, 1.034061e-07, 2.133243e-08, -2.641741e-08, 6.180585e-08, 
    -4.340427e-08, 4.290541e-08, 8.895836e-08, 1.603689e-08, -8.0056e-09, 
    8.128245e-08, 1.309816e-08, -5.704209e-09, -1.18024e-07, -2.343167e-08, 
    1.738486e-07, -1.401963e-07, -1.207563e-07, -9.297427e-09, 5.619313e-09, 
    1.11072e-09, -1.159904e-07, -7.950234e-08, -9.733458e-09, -3.116796e-09, 
    3.659358e-08, 1.192484e-08, -2.67984e-08, 8.733227e-08, -5.10008e-08, 
    8.674306e-11, 1.059104e-07, 1.00513e-07, -7.309019e-07, 1.067494e-07, 
    5.882839e-09, -1.547487e-07, -3.538594e-08, 5.627389e-08, 3.926115e-08, 
    1.119622e-07, -3.86683e-08, 1.920353e-08, 2.681645e-08, 4.253138e-08, 
    7.923018e-08, 8.194002e-08, 2.831325e-08, -6.205528e-08, 3.414858e-08, 
    1.011153e-08, 1.243706e-09, 1.873343e-08, -1.137528e-08, -2.150509e-07, 
    -2.683531e-07, 2.130055e-08, -1.030558e-07, -1.309559e-08, -8.581287e-08, 
    3.978244e-08, 3.039463e-08, 2.333491e-08, -6.50476e-08, -1.398338e-07, 
    2.220349e-07, -4.202379e-08, 9.81828e-09, 2.236548e-07, 7.314543e-08, 
    2.739656e-07, 7.349458e-08, -1.519788e-08, -1.154485e-07, 8.430606e-09, 
    -2.214938e-08, -6.992171e-08, -4.343858e-08, -9.51546e-09, 1.545004e-09, 
    -1.60253e-08, 3.041168e-08, -4.865797e-10, -4.897288e-08, -4.714639e-08, 
    -2.291517e-08, -7.724725e-08, 1.74964e-09, 5.291486e-08, -3.172681e-08, 
    -2.779734e-09, 5.400125e-13, -1.285002e-09, 1.072763e-09, 2.374372e-08,
  -8.506163e-09, 1.026592e-10, -2.702302e-08, 2.088211e-08, 4.346532e-08, 
    1.753403e-08, -4.150741e-08, 1.254432e-08, 4.523486e-09, 6.102789e-08, 
    7.996584e-08, 2.380738e-07, -5.004279e-08, -2.274504e-07, 6.626885e-08, 
    3.122195e-08, 2.930474e-08, 9.444784e-08, -1.4199e-08, -2.229095e-07, 
    -7.161054e-08, 1.177995e-07, -1.142949e-07, 2.346667e-08, 3.125862e-07, 
    2.108665e-07, 1.036143e-07, 2.194804e-08, -5.286404e-08, 9.871076e-08, 
    -3.86184e-08, 1.340574e-07, 4.935794e-08, 1.781666e-08, 1.834565e-09, 
    1.066804e-07, 3.561538e-08, -5.611753e-09, -1.224615e-07, -1.819008e-08, 
    1.095019e-07, -2.102462e-07, -5.536583e-08, -6.175618e-09, 1.740489e-08, 
    -9.158725e-09, -1.600312e-07, -6.348643e-08, -1.325118e-08, 
    -3.815884e-09, 3.720274e-08, 1.47337e-08, -2.830593e-08, 9.104622e-08, 
    -4.601746e-08, -2.176762e-09, 8.147765e-08, 3.357841e-08, -1.194793e-06, 
    8.518708e-08, 3.740058e-08, -3.805997e-08, 5.221489e-08, 3.679468e-08, 
    6.371944e-08, 5.362392e-08, -3.064054e-08, 1.114756e-08, 7.947051e-09, 
    3.526713e-08, 7.735969e-08, 1.118357e-07, 3.473372e-08, -4.075639e-08, 
    1.522297e-07, 1.115961e-08, 8.483312e-09, 1.466418e-08, -1.482484e-08, 
    -6.525318e-08, -2.841782e-07, 2.657439e-08, -1.188828e-07, -2.590127e-09, 
    -7.018673e-08, 4.21652e-08, 1.536902e-07, 1.427372e-08, -6.774862e-08, 
    -1.30176e-07, 2.055742e-08, -4.483134e-08, 1.96643e-08, 1.8943e-07, 
    2.187073e-08, 2.804248e-07, 5.025652e-08, 1.52678e-08, -8.632958e-08, 
    3.727338e-10, 6.687173e-09, -2.500035e-08, -4.270831e-08, -1.254736e-08, 
    5.287563e-08, 3.590117e-09, 3.114531e-08, -1.137539e-08, -5.414734e-08, 
    -4.935976e-08, -1.656497e-08, -6.273365e-08, -8.906568e-09, 4.627168e-09, 
    -3.724438e-08, -2.442562e-09, 9.890755e-12, -2.378378e-09, 1.146745e-09, 
    -2.269837e-08,
  -1.941402e-08, 3.182998e-08, -4.188706e-08, -1.730717e-08, 8.305659e-08, 
    6.472027e-08, -3.371446e-08, 4.395878e-08, -1.792267e-08, 2.242854e-08, 
    8.507055e-08, -1.258417e-08, -4.10152e-08, 8.280705e-08, -8.031617e-08, 
    3.965158e-08, 5.301042e-08, 1.110769e-07, 9.230493e-08, -1.49551e-07, 
    -2.093321e-08, -5.7264e-08, -4.416694e-08, 2.82534e-08, 7.375462e-08, 
    7.421403e-08, 8.62488e-08, 2.246628e-08, -7.072123e-08, 9.255433e-08, 
    -3.23169e-08, 5.433554e-08, 8.170554e-08, 7.239333e-08, 1.904942e-08, 
    1.839281e-07, 5.718813e-08, -4.390344e-09, -1.140804e-07, -3.262098e-08, 
    7.790288e-08, -9.859451e-08, -5.184091e-08, 1.987058e-09, -1.645896e-08, 
    -3.102656e-08, -1.244083e-07, -5.544229e-08, -2.773885e-08, 
    -4.178965e-09, 3.717514e-08, -5.526152e-08, -3.066156e-08, 9.190376e-08, 
    -3.275927e-08, -9.675603e-09, 5.341059e-08, 3.021572e-08, -1.190926e-06, 
    -8.07126e-08, 4.267685e-08, -6.84808e-08, 7.909597e-08, 6.280414e-09, 
    8.196196e-08, 3.510166e-08, 2.317978e-08, 2.170111e-09, 1.093446e-08, 
    3.242536e-08, 7.229227e-08, 1.263178e-07, 1.48238e-08, 7.025278e-10, 
    1.621054e-07, 1.69062e-08, 3.70494e-09, -1.068923e-08, -1.16615e-08, 
    4.380587e-08, -2.779061e-07, 1.790004e-08, -1.091464e-07, -2.625853e-08, 
    -2.226335e-08, -1.863822e-08, 1.157808e-07, 5.013987e-09, -7.337145e-08, 
    -9.802613e-08, 1.275947e-07, -2.964501e-08, 2.15957e-08, 1.573898e-07, 
    -4.233522e-08, 3.098228e-07, 2.672388e-08, 1.073539e-08, -5.33152e-08, 
    6.021613e-08, 1.178449e-08, -6.36098e-08, -3.886067e-08, -1.236979e-08, 
    -6.543871e-09, 2.535984e-08, 2.892477e-09, -2.61702e-08, -5.922385e-08, 
    -5.211831e-08, -1.403311e-08, -2.747078e-08, -1.263874e-08, 
    -3.087069e-08, -9.148778e-09, 1.899479e-10, 1.056165e-09, -2.66272e-09, 
    1.395129e-09, 1.626842e-08,
  -6.583207e-09, 6.067916e-08, -6.116016e-08, 7.949592e-08, 3.023751e-07, 
    1.273501e-07, -1.875952e-08, 1.538828e-07, -7.897654e-09, 4.795169e-08, 
    8.181303e-09, -1.148243e-08, 1.186476e-07, 2.086716e-08, -7.982914e-08, 
    4.75606e-08, 6.646752e-08, 4.65804e-08, 6.813747e-08, -4.159511e-08, 
    -8.934882e-08, -1.107601e-07, -3.710039e-08, -1.270201e-07, 3.73683e-09, 
    -1.721333e-07, 8.529167e-08, 1.532447e-08, -7.174464e-08, 4.842667e-08, 
    -1.454106e-08, 7.129796e-08, 9.831336e-08, 7.013563e-08, 5.127089e-08, 
    2.315869e-07, 6.945319e-08, -3.041777e-09, -9.213937e-08, -5.407177e-08, 
    1.233181e-07, -1.042332e-08, -7.061772e-08, 1.3774e-08, -7.943356e-09, 
    -4.58586e-08, -6.427666e-08, -3.929512e-08, -3.656556e-08, -5.220883e-09, 
    3.650641e-08, -1.214863e-07, -2.302601e-08, 8.526298e-08, -3.194883e-08, 
    1.086562e-09, 4.63462e-08, 4.63543e-08, -8.798281e-07, -3.732026e-08, 
    3.34723e-08, -8.758826e-08, -7.989513e-09, -4.67727e-09, 8.746436e-08, 
    4.177281e-08, 2.74278e-08, -2.494801e-09, 3.016424e-08, 3.38618e-08, 
    3.964095e-08, 1.076011e-07, 1.019947e-08, 7.001034e-08, 5.144221e-08, 
    2.05211e-08, -2.663114e-10, -5.969014e-09, 3.050815e-09, 1.075377e-07, 
    -2.546411e-07, 7.239402e-09, -1.130866e-07, -7.079512e-08, 1.347524e-08, 
    -7.368328e-09, 9.133436e-08, -3.286743e-09, -6.253475e-08, -2.423513e-08, 
    -4.152577e-08, -2.939515e-08, 1.839203e-08, 9.274081e-08, 4.87193e-08, 
    3.236374e-07, 7.814594e-09, 5.308556e-08, -3.705469e-08, 4.568991e-08, 
    8.486376e-08, 1.098786e-08, -3.322634e-08, -9.254251e-09, -6.798069e-08, 
    1.213875e-07, -7.04182e-09, -3.86047e-08, -6.351121e-08, -5.515204e-08, 
    -1.286895e-08, -1.29333e-08, 5.064749e-11, 8.289476e-10, 4.524168e-10, 
    1.275623e-09, -5.896396e-09, -2.752117e-09, 1.569418e-09, 7.884086e-08,
  -5.467462e-08, -8.601114e-08, 4.065593e-07, 6.648504e-07, 6.247278e-07, 
    8.61337e-09, -6.368543e-08, 8.218421e-09, 8.675408e-08, 4.664855e-08, 
    -2.240427e-08, -5.846073e-08, 4.860954e-08, -1.165255e-07, -3.787636e-08, 
    3.753266e-08, 8.431535e-08, 1.941152e-08, 6.721937e-08, 1.712112e-08, 
    -1.154968e-07, -1.420631e-08, 3.418506e-08, 2.707816e-08, -1.727813e-09, 
    -2.020042e-07, 7.083406e-08, 1.344176e-08, -5.982588e-08, -8.483084e-09, 
    1.559101e-09, 1.050686e-07, 1.692749e-07, 2.12319e-07, 7.41702e-08, 
    8.839208e-08, 7.309666e-08, -2.686662e-09, -6.96507e-08, -6.381458e-08, 
    1.388735e-07, 5.208506e-08, -9.087253e-08, 2.398284e-08, -1.592116e-08, 
    -2.477543e-08, -3.388601e-08, -2.603997e-08, -3.911898e-08, 
    -4.928047e-09, 3.543229e-08, -8.175959e-08, -1.462636e-08, 7.070455e-08, 
    -3.163727e-08, 1.047738e-09, 5.108859e-08, 4.447275e-08, -4.203459e-07, 
    -4.702208e-08, -9.39466e-08, -2.394131e-08, -2.671288e-08, 3.472337e-09, 
    9.197058e-08, 3.78775e-08, 2.488889e-08, -8.133497e-09, -2.6865e-08, 
    3.324101e-08, -1.379817e-08, 3.161392e-08, -3.042703e-08, -8.975451e-08, 
    1.344669e-08, 2.797094e-08, 1.017008e-08, 1.632372e-09, 6.542968e-09, 
    5.693437e-09, -2.090893e-07, -1.470117e-08, -1.224287e-07, 2.378704e-08, 
    1.245961e-07, 1.047167e-07, 2.886929e-08, -2.125296e-08, -2.871921e-08, 
    -1.746764e-08, -4.837625e-08, -2.079266e-08, 1.369506e-08, 6.362717e-08, 
    1.131184e-08, 3.178124e-07, -4.033413e-08, -2.866534e-08, -4.098399e-08, 
    1.244007e-08, 1.198823e-07, 1.037143e-07, -2.721058e-08, -7.659182e-09, 
    -5.668551e-08, 1.205e-07, -3.771561e-09, -5.020263e-08, -6.813718e-08, 
    -5.868742e-08, -1.183616e-08, -9.23751e-09, 3.502237e-09, 2.119805e-09, 
    2.274192e-09, 1.959643e-09, -4.034149e-09, -3.551669e-09, 1.434657e-09, 
    1.335138e-08,
  -1.760796e-07, -9.926994e-07, 1.671646e-07, 3.098522e-07, 1.893564e-07, 
    -3.659574e-08, -4.997122e-08, -4.473515e-08, -1.359359e-08, -1.73174e-08, 
    -1.799123e-08, -1.055549e-07, 2.070635e-09, -5.87649e-08, -4.269452e-09, 
    1.131104e-09, 9.959144e-08, -3.328694e-09, -2.291966e-08, 2.743076e-08, 
    1.104542e-08, -2.217331e-08, 2.411986e-08, -1.370273e-08, -4.970218e-09, 
    -1.179328e-07, 1.061579e-08, 1.073118e-08, -4.430757e-08, 2.074347e-08, 
    9.493419e-10, 6.407237e-08, 7.915838e-08, 5.71793e-07, 2.935613e-07, 
    -3.352937e-08, 7.294356e-08, -2.173806e-09, -3.902557e-08, -6.829905e-08, 
    1.411059e-07, 2.067935e-08, -8.897268e-08, 2.420289e-08, -6.249195e-09, 
    7.294074e-08, -1.775749e-08, -5.237951e-09, 1.594896e-08, -2.182432e-09, 
    3.406716e-08, 7.846268e-09, -7.079314e-09, 5.626331e-08, -2.438231e-08, 
    -1.444619e-09, 4.16091e-08, 5.308005e-08, -2.829799e-07, 5.547388e-08, 
    -3.774113e-08, -4.261216e-08, 2.374922e-07, 8.486071e-08, 1.071362e-07, 
    2.640144e-08, -7.116228e-10, -2.523791e-09, -2.540372e-08, 3.679526e-08, 
    -6.103676e-09, -2.347923e-08, -6.416366e-08, -7.036391e-08, 
    -3.636202e-08, 1.087375e-08, 1.524516e-08, 3.17533e-09, 6.959755e-09, 
    -1.888208e-08, -1.734135e-07, -8.466716e-09, -1.372765e-07, 4.558029e-08, 
    8.065268e-08, 9.544777e-08, -5.502335e-08, -6.104511e-08, 3.703983e-08, 
    -3.094357e-08, -4.099564e-08, -3.358597e-08, 1.258479e-08, 7.101778e-08, 
    -1.047732e-08, 3.170192e-07, -9.833487e-08, -5.37737e-08, -3.525184e-08, 
    1.403999e-09, 1.169669e-07, 1.212223e-08, 1.524024e-07, -6.258141e-09, 
    -5.163889e-08, 5.575833e-08, 7.298297e-09, -6.067904e-08, -7.335922e-08, 
    -6.264389e-08, -1.098039e-08, -7.600704e-09, 4.686569e-09, 2.575064e-09, 
    2.788227e-09, 2.394267e-09, -3.078682e-09, -3.324313e-09, 1.114167e-09, 
    -3.271845e-08,
  -2.381113e-07, -9.041013e-07, -9.731474e-08, -4.264842e-08, 5.058496e-10, 
    7.60835e-08, -1.067798e-08, 2.00659e-08, 1.308791e-08, -2.797861e-08, 
    -7.794739e-08, -2.43327e-07, -1.702773e-08, -3.293792e-09, 1.256238e-07, 
    -4.743921e-10, 1.203741e-07, -2.106373e-08, 7.381303e-09, -7.772206e-08, 
    3.960969e-08, -4.969309e-09, 2.290579e-08, 3.729497e-10, -9.672988e-09, 
    -1.245942e-07, -1.31898e-07, 7.721894e-09, -3.076553e-08, 2.749363e-08, 
    -2.280757e-08, 1.277803e-07, -3.007852e-08, 3.153586e-07, 2.947809e-07, 
    -5.913222e-08, 7.064924e-08, -1.413113e-09, -7.579445e-09, -7.159805e-08, 
    3.576446e-08, 1.66454e-08, -3.470117e-08, 1.444302e-08, -1.300651e-08, 
    6.205352e-08, -5.935703e-09, 1.289578e-08, 8.771232e-08, 1.495003e-09, 
    3.240743e-08, 1.710216e-07, -2.882996e-09, 4.505933e-08, -2.269444e-08, 
    -3.31454e-10, 2.749795e-08, 8.256266e-08, -3.44742e-07, 4.929265e-08, 
    -3.733504e-08, 3.099348e-08, -6.37823e-09, 1.927473e-08, 1.219714e-07, 
    3.289358e-09, -1.416396e-08, 2.310099e-08, 1.057987e-08, 2.941186e-08, 
    -4.204082e-09, -2.664314e-08, -7.948194e-08, -7.413411e-08, 
    -5.313491e-08, -6.228504e-09, 6.476102e-08, 7.672185e-09, 3.564166e-08, 
    -8.423973e-08, -1.594581e-07, 2.74627e-08, -1.490716e-07, 2.571207e-07, 
    -2.267001e-08, 1.041697e-07, -8.875605e-08, -9.988361e-08, -2.273886e-08, 
    -4.383708e-08, 1.874304e-08, -4.49062e-08, 3.155085e-08, 4.867106e-08, 
    -1.177415e-08, 3.256313e-07, -1.286909e-07, -1.768257e-08, -1.469118e-09, 
    6.829589e-09, -1.356801e-08, -3.885013e-09, 7.336407e-08, -7.317098e-09, 
    -3.035353e-08, -6.628682e-09, 1.613643e-08, -7.160321e-08, -7.912371e-08, 
    -6.724844e-08, -1.09506e-08, -6.798871e-09, 5.322306e-09, 3.028788e-09, 
    2.976151e-09, 3.004516e-09, -1.05878e-09, -2.264237e-09, 3.786269e-10, 
    1.325822e-08,
  -1.930845e-07, 3.398395e-08, -1.0592e-07, -1.094281e-08, -4.449646e-08, 
    1.38524e-08, 1.345109e-08, 3.240757e-09, 7.125323e-09, 1.980015e-08, 
    -8.800691e-08, -6.204992e-07, -8.828351e-09, -3.634568e-10, 
    -4.794174e-10, 1.372379e-08, 1.210167e-07, 2.678365e-08, 4.679939e-08, 
    4.539311e-08, -1.03413e-08, 2.293632e-09, 2.471756e-08, 6.808136e-09, 
    -8.76696e-09, -6.814491e-08, -2.228387e-08, -7.357812e-10, -2.066565e-08, 
    -3.912191e-09, -7.356402e-08, 3.077749e-07, -4.768094e-08, 1.764723e-07, 
    -8.141615e-08, 9.792313e-08, 6.267901e-08, -1.168985e-10, 1.922933e-08, 
    -6.336804e-08, 4.550233e-08, 1.535682e-08, -1.799663e-08, 1.109926e-08, 
    -6.538357e-09, 5.004199e-08, -1.113278e-09, 3.086527e-08, 7.34731e-08, 
    3.933799e-09, 3.173677e-08, 4.86101e-08, -1.125284e-09, 3.334933e-08, 
    -2.19034e-08, -5.352376e-09, 9.98989e-09, 7.266421e-08, -4.256259e-07, 
    -9.284221e-09, -1.882768e-08, 3.566242e-08, -2.536876e-08, -2.346314e-09, 
    1.300458e-07, -3.026287e-08, -3.842501e-08, -1.207673e-08, -8.127131e-09, 
    2.16661e-08, -1.008789e-08, -2.516947e-08, -3.584307e-08, 1.232047e-08, 
    -6.111802e-08, -1.197952e-08, 3.300299e-08, -2.535756e-09, 1.55517e-08, 
    -3.085233e-08, -1.67446e-07, 7.700769e-08, -1.479921e-07, 3.777359e-09, 
    -1.012756e-08, 7.93367e-08, -1.435079e-07, -6.81141e-08, -5.965919e-08, 
    -5.03673e-08, -1.983494e-09, -2.556076e-08, -7.72522e-09, 4.442696e-08, 
    -2.659442e-08, 3.116636e-07, -1.217594e-07, 1.030294e-07, 1.282535e-08, 
    9.721679e-09, -6.590153e-08, -1.001128e-08, 1.096979e-08, -6.858173e-09, 
    -9.130133e-08, -4.595734e-08, 1.923604e-08, -8.68389e-08, -8.666905e-08, 
    -7.23528e-08, -1.118531e-08, -6.377491e-09, 6.463893e-09, 3.306127e-09, 
    3.904006e-09, 2.855063e-09, 3.580737e-09, -1.302162e-09, 6.343015e-11, 
    1.487172e-08,
  -1.41183e-07, 3.502743e-08, -1.006973e-07, -2.051496e-08, -1.808365e-08, 
    4.946912e-09, 4.19692e-09, -4.911328e-09, 4.494439e-09, 3.412481e-09, 
    -4.959986e-09, -3.597422e-07, -1.255302e-08, 2.952049e-09, -1.491372e-08, 
    9.894631e-09, 1.016909e-07, 1.96722e-08, 4.299451e-08, 7.955106e-08, 
    -5.602772e-09, 3.61814e-09, 2.658265e-08, 9.371149e-09, -1.011466e-08, 
    1.584073e-08, 6.699469e-08, -1.10785e-08, -1.790846e-08, 4.008604e-08, 
    -1.000471e-07, 1.91086e-07, -1.072218e-07, 9.455908e-08, -7.960438e-08, 
    1.635331e-07, 5.136475e-08, 6.835421e-12, 1.484028e-08, -5.751871e-08, 
    -4.212936e-08, 1.497784e-08, -1.803954e-08, 3.358245e-09, -9.511666e-09, 
    1.248048e-08, -9.945325e-10, 4.892888e-08, 1.997958e-08, 5.479038e-09, 
    3.147977e-08, -3.626855e-08, -1.37095e-09, 2.307657e-08, -2.127507e-08, 
    -3.255252e-09, -5.58083e-09, 6.749113e-08, -4.728487e-07, 2.948994e-09, 
    -1.231405e-08, 3.590861e-08, -3.006727e-08, -8.74444e-09, 1.205286e-07, 
    -3.561337e-08, -6.093723e-08, -6.313184e-08, 2.772543e-08, -1.71828e-08, 
    2.550547e-08, -2.387839e-08, 1.365492e-07, 2.411736e-08, -6.543811e-08, 
    7.103324e-09, 4.604701e-09, -1.595311e-10, 1.451779e-08, 5.247472e-08, 
    -1.44255e-07, 4.010898e-08, -1.530124e-07, -2.049109e-08, -1.842881e-08, 
    1.940995e-07, 5.163469e-08, 3.452595e-08, -4.901678e-08, -5.647934e-08, 
    1.62612e-09, -9.646158e-09, -4.08474e-09, 5.818726e-08, 1.354553e-07, 
    2.720161e-07, -1.028971e-07, 8.070214e-08, -6.082757e-09, -1.847908e-08, 
    -1.142155e-09, -1.205175e-08, -4.838079e-08, -6.582944e-09, 1.686175e-08, 
    -6.964405e-08, 2.568703e-08, -9.356467e-08, -8.823116e-08, -7.8406e-08, 
    -1.190875e-08, -6.343782e-09, 7.91232e-09, 3.550838e-09, 1.543356e-09, 
    2.599745e-09, 6.097665e-09, -1.167578e-09, 8.773355e-10, 1.772122e-08,
  -2.108049e-07, 1.955419e-08, -5.216583e-08, -4.157431e-08, -1.096322e-08, 
    1.450019e-09, 5.098855e-11, -8.274299e-09, 4.19692e-09, 4.877677e-09, 
    3.606431e-09, -2.239546e-07, -1.320831e-08, 8.497466e-09, -1.809275e-08, 
    -9.602321e-09, 7.97671e-08, -1.988809e-08, 4.813973e-08, 8.486137e-08, 
    -6.731796e-09, 7.056144e-09, 2.800249e-08, 9.763255e-09, -1.402253e-08, 
    2.017015e-08, 8.557896e-08, -7.457692e-08, -2.108567e-08, 4.721284e-08, 
    -1.352323e-07, 1.662038e-07, -9.138392e-08, 9.966612e-08, -7.828766e-08, 
    2.018301e-07, 3.948456e-08, -9.075052e-11, -2.833229e-08, -5.479961e-08, 
    -5.760384e-08, 1.567111e-08, -3.42194e-08, -2.841954e-08, 4.682363e-09, 
    -5.720437e-09, -3.196021e-09, 6.206102e-08, -4.348748e-08, 6.16636e-09, 
    3.154949e-08, -4.579914e-08, -2.181229e-09, 1.632467e-08, -2.084551e-08, 
    -5.482718e-09, -2.245605e-08, 5.601311e-08, -4.872941e-07, 9.389396e-10, 
    -1.307802e-08, 3.407337e-08, -3.1561e-08, 2.136486e-08, 9.297125e-08, 
    4.78056e-08, -6.047998e-08, 4.849568e-08, 9.078423e-08, -2.565997e-08, 
    2.703047e-08, -2.296741e-08, 1.579684e-08, 2.588132e-08, -6.800762e-08, 
    -5.64313e-09, 3.722562e-09, -8.735014e-09, -5.569609e-09, 6.749644e-09, 
    -1.341734e-07, 3.067351e-08, -1.562228e-07, -2.624705e-08, -2.052974e-08, 
    3.39071e-10, 8.593162e-08, 3.466454e-08, -5.203515e-08, -6.193608e-08, 
    3.447951e-09, -5.274103e-09, -5.799279e-09, 6.390108e-08, 9.381148e-08, 
    2.405891e-07, -9.392178e-08, 1.252886e-09, -2.590326e-08, -1.488864e-08, 
    3.03167e-08, -1.379532e-08, -7.929498e-08, -6.693327e-09, 1.540258e-08, 
    -1.075122e-07, 3.691963e-08, -8.817773e-08, -7.661123e-08, -8.038609e-08, 
    -1.310372e-08, -6.419612e-09, 9.013149e-09, 3.448633e-09, -2.718821e-10, 
    2.778404e-09, 2.543658e-09, -2.976833e-09, 1.061863e-09, 1.836207e-08,
  -1.151836e-07, 1.192461e-08, -4.275762e-08, -4.729986e-08, -6.316441e-09, 
    -2.262368e-10, -5.337597e-09, -9.588121e-09, 1.385843e-09, 3.046807e-11, 
    2.551224e-08, -1.442995e-07, -1.279864e-08, 7.364406e-09, -1.786862e-08, 
    -4.292667e-08, 6.041359e-08, -2.274408e-08, 4.935848e-08, 9.198288e-08, 
    -7.524477e-09, 8.185907e-09, 2.909019e-08, 1.061585e-08, -1.666513e-08, 
    2.233946e-08, 9.801943e-08, -8.679081e-08, -4.497019e-08, 4.927847e-08, 
    -1.37381e-07, 8.777897e-08, -1.830676e-08, 1.055034e-07, -7.688959e-08, 
    2.277172e-07, 2.750382e-08, -2.660272e-10, -4.118215e-08, -4.338585e-08, 
    -8.023909e-08, 1.633612e-08, -7.399962e-08, -1.55011e-08, 3.288801e-08, 
    8.089273e-09, -6.702635e-09, 6.57576e-08, -5.595439e-08, 6.734894e-09, 
    3.178431e-08, -4.987578e-08, -3.570745e-09, 1.172511e-08, -2.048756e-08, 
    -5.212428e-09, -4.241656e-08, 6.296252e-08, -4.913722e-07, 3.382411e-09, 
    -1.233116e-08, 3.231253e-08, -3.183914e-08, 1.96635e-08, 7.452654e-08, 
    3.188893e-08, -3.921468e-08, 5.502284e-08, 5.39917e-08, 1.082412e-08, 
    5.607626e-08, -2.30807e-08, -5.896027e-08, 2.603451e-08, -6.967377e-08, 
    -1.452781e-08, 3.546603e-09, -1.215739e-08, -1.762104e-08, -2.481784e-09, 
    -1.076762e-07, 3.44275e-08, -1.568174e-07, -2.849652e-08, -2.108072e-08, 
    -3.286459e-09, 8.403936e-08, 3.331388e-08, -6.009614e-08, -6.434789e-08, 
    4.707317e-09, -3.419881e-09, -6.174616e-09, 7.960688e-08, -9.846508e-08, 
    2.19337e-07, -8.932048e-08, -1.939088e-08, -3.732839e-08, -1.224503e-08, 
    3.625587e-08, -1.48714e-08, -8.664152e-08, -6.641244e-09, 1.974308e-08, 
    -1.122332e-07, 4.917501e-08, -8.44293e-08, -6.974892e-08, -6.9105e-08, 
    -1.19046e-08, -6.35373e-09, 9.200676e-09, 3.383093e-09, -2.678462e-09, 
    5.356878e-09, 1.774396e-09, -3.880551e-09, 4.753957e-10, 1.583362e-08,
  -6.581996e-08, 8.461427e-09, -3.732492e-08, -4.515636e-08, -3.377806e-09, 
    -1.173419e-09, -6.935636e-09, -7.432561e-09, 1.292221e-09, -3.143612e-09, 
    3.061103e-08, -5.584963e-08, -1.591769e-08, 5.475215e-09, -2.163512e-08, 
    -7.472254e-08, 4.712345e-08, -2.35313e-08, 5.02947e-08, 9.733475e-08, 
    -8.152426e-09, 7.696087e-09, 2.92211e-08, 1.159304e-08, -1.659549e-08, 
    2.17828e-08, 7.618263e-08, 9.111676e-08, -5.607916e-08, 7.411944e-08, 
    -1.203913e-07, 6.135355e-08, -2.71054e-07, 1.128541e-07, -7.552291e-08, 
    2.919816e-07, 1.707092e-08, 3.222027e-10, -4.682994e-08, -4.120768e-08, 
    -1.092926e-07, 1.454254e-08, -6.805186e-08, -8.284742e-09, 5.820056e-08, 
    2.607504e-08, -1.052229e-08, 6.832386e-08, -7.21973e-08, 7.287866e-09, 
    3.207408e-08, -5.251746e-08, -5.326217e-09, 9.091821e-09, -2.021125e-08, 
    -1.307797e-09, -5.30826e-08, 6.47459e-08, -4.858416e-07, 1.466603e-09, 
    -1.214488e-08, 3.288295e-08, -3.157373e-08, 2.659973e-08, 6.573949e-08, 
    1.080315e-08, -3.690104e-09, 4.089674e-08, 3.435474e-08, 1.824998e-08, 
    -1.039666e-10, -2.454891e-08, -5.612452e-08, 2.573501e-08, -7.048118e-08, 
    -1.672964e-08, 3.960579e-09, -1.238539e-08, -1.123437e-08, -7.127653e-09, 
    -9.564377e-08, 3.590671e-08, -1.559021e-07, -2.963731e-08, -2.104963e-08, 
    -8.425843e-09, 6.425461e-08, 3.178178e-08, -6.200685e-08, -6.681597e-08, 
    5.849472e-09, -3.782532e-09, -6.347562e-09, 8.935741e-08, -1.072725e-07, 
    1.867151e-07, -6.963859e-08, -1.670418e-08, -5.07485e-08, -1.007021e-08, 
    4.244481e-08, -1.254095e-08, -9.192015e-08, -6.031023e-09, 2.875885e-08, 
    -1.129582e-07, 6.945828e-08, -8.875423e-08, -6.804413e-08, -6.048441e-08, 
    -8.323752e-09, -5.544791e-09, 7.662322e-09, 3.308116e-09, -8.127188e-09, 
    1.15823e-09, 7.853544e-09, -1.047065e-08, 1.644771e-09, 1.891732e-08,
  -5.655011e-08, 7.484346e-09, -3.481296e-08, -4.184346e-08, -1.43973e-09, 
    -1.505441e-09, -6.396817e-09, -6.09225e-09, 7.148628e-10, -6.080541e-09, 
    3.763478e-08, -2.199977e-08, -1.511489e-08, 5.004949e-09, -2.584704e-08, 
    -8.159435e-08, 4.034166e-08, -2.375123e-08, 5.022252e-08, 1.014437e-07, 
    -8.500251e-09, 7.574045e-09, 2.836782e-08, 1.265448e-08, -1.592616e-08, 
    2.399781e-08, 9.670021e-08, 1.015344e-07, -4.811932e-08, 8.442328e-08, 
    -1.056735e-07, -1.077547e-08, -3.007376e-07, 1.130005e-07, -7.434073e-08, 
    3.082846e-07, 8.985467e-09, -7.196377e-11, -4.57643e-08, -4.019513e-08, 
    -1.294676e-07, 1.399974e-08, -6.860068e-08, -5.004775e-09, 3.537559e-08, 
    4.510787e-08, -1.497483e-08, 6.709536e-08, -7.86956e-08, 7.135476e-09, 
    3.272967e-08, -5.440791e-08, -6.783318e-09, 8.616894e-09, -2.003112e-08, 
    -5.230163e-10, -5.827394e-08, 6.040534e-08, -4.754038e-07, -4.976926e-10, 
    -1.242563e-08, 3.477646e-08, -3.087939e-08, 2.539407e-08, 5.948159e-08, 
    -3.522814e-09, -1.100518e-07, 2.543982e-08, 2.567469e-08, -5.968786e-09, 
    -4.744152e-09, -1.904584e-08, -5.775848e-08, 2.53076e-08, -7.051207e-08, 
    -1.242529e-08, 4.274369e-09, -1.17424e-08, -1.335895e-08, -1.058208e-08, 
    -9.674818e-08, 3.883154e-08, -1.546186e-07, -3.033904e-08, -2.064553e-08, 
    -1.139847e-08, 4.940057e-08, 3.04542e-08, -6.168862e-08, -6.808261e-08, 
    4.65684e-09, -3.438821e-09, -6.43152e-09, 9.548647e-08, -1.521498e-07, 
    1.606873e-07, -6.049902e-08, -3.949015e-08, -5.382026e-08, -7.43437e-09, 
    4.564799e-08, -1.216137e-08, -9.428239e-08, -4.589083e-09, 3.198704e-08, 
    -1.128157e-07, 2.255759e-07, -9.583539e-08, -6.861444e-08, -5.870311e-08, 
    -5.142738e-09, -4.100116e-09, 8.306984e-09, 3.332957e-09, -1.510682e-08, 
    -8.304027e-10, 1.390394e-08, -9.518821e-10, 7.102187e-09, 2.265415e-08,
  -4.26794e-08, 5.707989e-09, -3.578225e-08, -4.173785e-08, -7.580638e-10, 
    -1.868102e-09, -2.816023e-09, -7.054496e-09, 1.10299e-09, -5.190259e-09, 
    3.724972e-08, 2.486104e-09, -1.46772e-08, 4.555886e-09, -2.915522e-08, 
    -5.488246e-08, 3.712705e-08, -2.391607e-08, 4.989636e-08, 1.046615e-07, 
    -8.783672e-09, 7.239123e-09, 2.650813e-08, 1.305284e-08, -1.478907e-08, 
    2.421848e-08, 1.078133e-07, 8.217557e-08, -4.350272e-08, 8.923098e-08, 
    -9.05527e-08, -3.090736e-08, -2.84914e-07, 1.218925e-07, -7.291692e-08, 
    3.337423e-07, 2.604452e-09, -1.094918e-09, -4.893582e-08, -4.056239e-08, 
    -1.645107e-07, 1.394847e-08, -6.84463e-08, 1.390333e-09, 2.957495e-08, 
    5.982156e-08, -1.989395e-08, 6.482094e-08, -8.460339e-08, 6.456318e-09, 
    3.414479e-08, -5.565812e-08, -8.033293e-09, 8.741154e-09, -1.989325e-08, 
    8.965344e-10, -6.430673e-08, 5.651884e-08, -4.605228e-07, -2.438696e-09, 
    -1.305261e-08, 3.718151e-08, -2.980141e-08, 2.440902e-08, 5.494663e-08, 
    2.183651e-08, -1.376752e-07, 4.085837e-08, 2.899947e-08, -1.12575e-08, 
    -7.674998e-09, 6.768232e-09, -6.185883e-08, 2.442084e-08, -6.985954e-08, 
    -1.610238e-08, 4.048616e-09, -1.125602e-08, -1.484266e-08, -1.296962e-08, 
    -1.020215e-07, 4.003241e-08, -1.535722e-07, -3.011291e-08, -2.050069e-08, 
    -1.298122e-08, 3.986906e-08, 2.875527e-08, -6.045347e-08, -6.853486e-08, 
    4.923095e-09, -8.890755e-10, -6.481059e-09, 1.03482e-07, -1.856208e-07, 
    1.595273e-07, -5.935749e-08, -6.731852e-09, -5.443667e-08, -7.07487e-09, 
    4.781009e-08, -1.230461e-08, -9.487296e-08, -5.065857e-09, 3.338778e-08, 
    -1.122457e-07, 5.940547e-08, -1.003918e-07, -6.910341e-08, -6.038999e-08, 
    -5.972879e-09, -3.92015e-09, 7.915332e-09, 2.972911e-09, -2.149864e-08, 
    3.383316e-11, 2.374239e-08, -3.830003e-09, 3.394902e-09, 2.300226e-08,
  -4.277518e-08, 4.059473e-09, -3.680208e-08, -4.26549e-08, 1.957119e-10, 
    -2.490026e-09, -4.379785e-10, -9.019288e-09, -1.193712e-12, 
    -5.321965e-09, 3.602344e-08, 1.757115e-08, -1.313566e-08, 4.360288e-09, 
    -2.860935e-08, 2.412943e-08, 3.489691e-08, -2.384223e-08, 4.944204e-08, 
    1.065397e-07, -8.481322e-09, 6.787047e-09, 2.467317e-08, 1.348343e-08, 
    -1.322093e-08, 2.195287e-08, 9.838794e-08, 7.845205e-08, -4.100826e-08, 
    9.155218e-08, -8.217359e-08, -4.603095e-08, -2.809539e-07, 1.262601e-07, 
    -7.101886e-08, 3.521031e-07, -3.512344e-09, -9.373196e-10, -3.971769e-08, 
    -3.614056e-08, -2.060345e-07, 1.369762e-08, -6.997709e-08, 4.56231e-09, 
    2.138239e-08, 7.24346e-08, -2.496978e-08, 6.196819e-08, -8.788798e-08, 
    7.379811e-09, 3.711682e-08, -5.612134e-08, -8.925565e-09, 1.309512e-08, 
    -1.981855e-08, 2.756622e-09, -6.844544e-08, 5.437763e-08, -4.398921e-07, 
    -2.988912e-09, -1.415134e-08, 3.954705e-08, -2.810231e-08, 2.337164e-08, 
    4.976063e-08, 3.617328e-08, -1.426106e-07, 4.627753e-08, 3.596432e-08, 
    -2.298594e-08, -7.246001e-09, -1.483915e-08, -5.642852e-08, 2.362657e-08, 
    -6.944289e-08, -1.500172e-08, 4.446974e-09, -1.097845e-08, -1.400152e-08, 
    -1.492668e-08, -9.703189e-08, 4.073608e-08, -1.549243e-07, -2.970802e-08, 
    -1.994096e-08, -1.31991e-08, 2.877044e-08, 2.622568e-08, -5.908762e-08, 
    -6.878662e-08, 7.360256e-09, -5.341114e-10, -6.518064e-09, 1.128895e-07, 
    -1.950535e-07, 1.385297e-07, -5.59624e-08, -1.302681e-09, -5.373596e-08, 
    -6.564424e-09, 5.026544e-08, -1.186923e-08, -9.270562e-08, -5.13937e-09, 
    3.519943e-08, -1.114141e-07, 4.204566e-08, -1.026588e-07, -6.947931e-08, 
    -6.132933e-08, -7.102756e-09, -4.572769e-09, 8.867744e-09, 1.526985e-09, 
    -2.550661e-08, 4.49188e-10, 2.049165e-08, 1.13871e-08, 2.615792e-10, 
    2.216979e-08,
  -4.315564e-08, -1.613785e-09, -3.917933e-08, -4.325523e-08, -7.486278e-10, 
    -3.2461e-09, -2.825118e-10, -7.698759e-09, -1.928697e-09, -5.823381e-09, 
    3.475213e-08, 2.551417e-08, -1.116075e-08, 3.856826e-09, -2.684635e-08, 
    5.877669e-08, 3.000646e-08, -2.311856e-08, 4.845657e-08, 1.030816e-07, 
    -7.263338e-09, 6.60259e-09, 2.339732e-08, 1.455339e-08, -1.20807e-08, 
    1.832984e-08, 1.057202e-07, 7.555684e-08, -3.967841e-08, 9.073494e-08, 
    -8.864106e-08, -5.150753e-08, -2.514201e-07, 1.230557e-07, -6.682751e-08, 
    3.760919e-07, -7.520339e-09, -1.450246e-09, -3.074331e-08, -4.325695e-08, 
    -2.86071e-07, 1.340879e-08, -6.349285e-08, 3.735014e-09, 2.105264e-08, 
    8.582572e-08, -3.00181e-08, 5.824285e-08, -9.305502e-08, 1.2491e-08, 
    4.470832e-08, -5.495883e-08, -9.559745e-09, 1.710894e-08, -1.988146e-08, 
    6.533128e-09, -6.896619e-08, 4.917204e-08, -4.061691e-07, -2.846321e-09, 
    -1.615729e-08, 3.989442e-08, -2.438958e-08, 2.243662e-08, 3.644334e-08, 
    4.342098e-08, -1.480076e-07, 4.429114e-08, 3.515731e-08, -2.595027e-08, 
    -2.940055e-09, -8.220798e-08, -5.957588e-08, 2.164086e-08, -6.678547e-08, 
    -1.50975e-08, 3.311612e-09, -9.856819e-09, -1.296804e-08, -1.700175e-08, 
    -8.820336e-08, 4.006461e-08, -1.503115e-07, -2.846366e-08, -1.916339e-08, 
    -1.108572e-08, 3.175944e-08, 2.095169e-08, -5.645416e-08, -6.895743e-08, 
    1.158207e-08, -6.379892e-10, -6.43422e-09, 1.148859e-07, -1.893058e-07, 
    6.675609e-08, -4.532096e-08, -2.960292e-09, -5.093591e-08, -6.859977e-09, 
    5.396817e-08, -9.62855e-09, -8.819787e-08, -4.895767e-09, 3.285993e-08, 
    -1.097038e-07, 3.584967e-08, -1.039294e-07, -6.981679e-08, -6.175298e-08, 
    -7.501171e-09, -4.779508e-09, 7.841322e-09, 9.856763e-09, -2.815966e-08, 
    2.362867e-10, 2.000056e-08, 5.480487e-10, 1.738985e-08, 2.00788e-08,
  2.43038e-13, -3.179147e-14, 5.161955e-14, 2.88763e-13, 2.70313e-13, 
    -4.506314e-14, -2.673842e-13, -5.276609e-13, -6.719638e-13, 
    -9.190223e-14, 4.55141e-13, 6.754126e-14, -1.263933e-13, -1.300225e-13, 
    1.63595e-13, -4.279546e-15, 2.724128e-13, -3.820351e-13, -2.819886e-13, 
    7.264306e-14, -3.702321e-13, -1.125392e-12, -5.422298e-13, 5.231999e-13, 
    -9.190737e-13, -6.810714e-13, -2.214376e-13, 1.633488e-13, 4.647401e-14, 
    3.275981e-14, -7.577295e-14, -1.5784e-13, -2.513782e-13, -7.343705e-14, 
    -1.884914e-13, -1.816058e-14, -1.203637e-13, -2.089219e-12, 4.790055e-13, 
    1.324197e-12, -5.321097e-13, 9.657971e-14, 1.832127e-13, 4.296982e-13, 
    1.441858e-13, 1.436488e-13, 1.764968e-13, 2.084393e-12, 3.034858e-13, 
    -4.438515e-13, -1.463551e-12, -4.8899e-13, 4.364867e-12, 1.575516e-12, 
    4.253009e-14, -5.701016e-13, 2.138129e-13, 9.808633e-13, 2.332568e-13, 
    -1.288745e-12, 1.03121e-12, 1.222306e-13, 2.998588e-13, -2.652104e-13, 
    -1.405289e-12, -5.851374e-14, -1.815138e-13, 3.024125e-13, 1.784024e-13, 
    6.727378e-14, -2.186782e-14, 1.150922e-14, 1.07266e-13, -1.104991e-13, 
    -5.371027e-13, 4.794054e-15, 1.153576e-12, 1.183344e-13, -2.641297e-12, 
    -9.921172e-13, -8.597827e-13, -1.998247e-12, -7.96355e-14, -6.421713e-13, 
    9.953017e-15, 2.92454e-13, 9.768119e-15, 8.169847e-13, 8.725031e-13, 
    3.55719e-12, -3.367192e-13, 1.948605e-13, -1.280729e-12, -1.139035e-12, 
    3.668206e-13, 2.984751e-13, 2.45916e-14, -1.3661e-13, 5.799761e-13, 
    5.027402e-13, -4.530804e-12, -4.07714e-13, 4.407241e-14, 3.182822e-13, 
    -7.368216e-14, 3.571803e-14, -1.267712e-13, -4.233028e-14, 2.570103e-14, 
    1.889354e-14, 9.422553e-14, 1.099384e-14, 1.468686e-13, 1.520591e-13, 
    6.478788e-13, -3.039714e-12, -1.020711e-13, 1.639399e-13, 1.765302e-13, 
    -3.191784e-13,
  8.60768e-14, 1.501958e-13, 1.292105e-13, 7.258163e-14, -9.548293e-14, 
    -1.365489e-13, -1.553135e-13, -1.185373e-13, -2.007038e-13, 
    -8.156514e-14, -6.381465e-15, -1.372055e-13, -3.942479e-13, 
    -3.196705e-13, -1.591899e-13, 1.395362e-13, 1.852465e-13, -2.956358e-13, 
    -7.197999e-13, -4.959622e-13, -4.420953e-13, -1.279888e-12, 
    -1.785692e-12, -6.617315e-14, 1.536443e-13, 1.892047e-13, 3.291068e-13, 
    3.340186e-13, 2.300478e-13, -6.214914e-14, -1.79769e-14, 3.148332e-14, 
    -1.163325e-13, 5.754407e-14, 1.782378e-13, 8.952251e-14, -2.066213e-12, 
    -7.310303e-13, 1.632132e-13, 2.252404e-13, -1.693243e-13, 1.09227e-13, 
    -7.583212e-13, 4.633286e-13, 7.728739e-14, 3.610959e-13, -4.424759e-13, 
    8.134456e-13, 1.620346e-13, 8.131074e-13, 3.477512e-14, -4.540057e-13, 
    1.559165e-12, -5.41596e-12, 3.561804e-13, -4.737456e-13, -3.243289e-13, 
    -6.336826e-13, 1.13292e-12, 3.188359e-12, 6.826936e-13, 1.715355e-13, 
    1.222919e-13, 1.586655e-13, 7.462129e-14, -6.645791e-13, -4.358717e-13, 
    -3.464582e-13, -2.332841e-14, 2.978286e-14, -7.657082e-13, 3.58414e-13, 
    8.229483e-13, 4.633117e-13, 9.918158e-13, -2.990951e-13, 3.377587e-13, 
    3.323277e-13, -4.286615e-12, 1.148974e-12, 5.179403e-13, 7.491847e-13, 
    -4.444547e-13, 4.803665e-13, 8.730238e-14, 1.203558e-12, -5.539172e-13, 
    -4.3115e-13, 7.092522e-14, 1.036807e-12, -1.226836e-14, -2.383364e-13, 
    4.97711e-13, 9.176693e-13, -2.231441e-13, 3.185216e-13, 1.701382e-13, 
    1.024712e-13, 4.846054e-13, 5.213317e-13, -3.95696e-13, 1.43967e-13, 
    -1.895443e-12, 1.670642e-13, -1.649685e-14, -5.108969e-13, 6.617736e-14, 
    -1.243585e-12, -9.343551e-13, -5.199788e-13, -6.306002e-13, 
    -1.140734e-13, 2.040675e-13, 2.146179e-13, 1.844573e-13, 7.958957e-13, 
    -1.924289e-13, -6.46139e-13, 7.648871e-14, -1.382586e-13,
  4.883594e-14, -9.832413e-14, -1.013217e-13, 5.77316e-15, 8.489043e-14, 
    1.98383e-13, 7.621681e-14, -3.376466e-14, -1.295491e-13, -1.858791e-13, 
    -4.395095e-14, 4.03011e-14, 5.193068e-14, 1.436351e-13, 9.105217e-14, 
    -1.115774e-14, 4.734477e-13, 4.049677e-13, 7.699015e-13, 1.017325e-12, 
    8.953532e-13, 8.366502e-13, 1.224937e-12, 2.936817e-13, 6.948053e-13, 
    5.152545e-13, 3.211598e-13, 2.815526e-13, 1.098149e-13, 1.527806e-13, 
    1.032646e-13, -7.713274e-14, 1.865313e-13, 5.24164e-14, 7.160939e-15, 
    9.17183e-14, -2.239439e-12, -1.113566e-12, -3.668177e-13, 7.31816e-13, 
    -3.162026e-13, -1.305345e-13, 5.938236e-13, 2.296414e-13, 6.307455e-14, 
    -1.359191e-13, -1.408963e-12, -5.503167e-13, -5.603268e-13, -3.01318e-13, 
    2.006416e-13, -2.897821e-13, 2.160036e-13, -8.99586e-12, 1.219153e-13, 
    1.244171e-12, -4.003048e-13, -1.184669e-12, 7.631423e-13, -2.547112e-13, 
    8.009843e-13, -2.723377e-13, 0, 5.413753e-13, 4.161699e-13, 
    -1.865869e-13, -1.139921e-13, -3.677614e-14, -3.033684e-14, 1.396105e-13, 
    6.728784e-13, 1.577211e-13, 5.043604e-13, 7.233519e-13, 3.787054e-13, 
    -2.828154e-12, -6.981568e-14, 4.780655e-13, 8.380137e-14, 5.17586e-13, 
    1.312249e-12, 7.213851e-13, -8.784085e-13, 6.093737e-13, 1.127307e-12, 
    1.563749e-13, 1.715891e-12, 6.404044e-13, 2.632781e-13, 1.021752e-13, 
    -3.944067e-14, -7.770173e-14, 2.202474e-13, -1.084709e-12, 9.710288e-14, 
    2.979103e-13, 1.616762e-14, -8.258672e-14, 5.96273e-13, 9.50004e-13, 
    -5.260792e-13, -1.584757e-14, 6.930567e-14, -4.666979e-13, -8.024414e-13, 
    -5.165451e-13, -6.447343e-13, -7.623485e-13, -1.419545e-12, 
    -8.607975e-13, 2.782635e-13, 6.256107e-14, 9.714451e-15, 1.481038e-13, 
    1.029912e-12, 1.695902e-12, 8.793138e-12, 4.296682e-12, -2.755704e-13, 
    -1.601802e-12,
  2.364775e-13, 2.066819e-13, 2.539358e-13, 2.638306e-13, 2.158829e-13, 
    1.242062e-13, 9.765799e-14, -9.003909e-14, -1.491862e-13, -1.999789e-13, 
    8.323897e-14, -2.510353e-13, -3.005513e-13, 1.333655e-13, -1.182804e-13, 
    2.741765e-13, 2.540343e-13, 8.276713e-14, 4.461986e-13, 6.522005e-13, 
    3.301109e-13, 4.278522e-13, 2.702838e-13, -2.99219e-13, -1.343176e-12, 
    -2.209621e-12, -9.54653e-14, 4.507644e-13, 1.863509e-13, 4.346246e-13, 
    3.524681e-13, -2.49939e-14, 3.937128e-14, 4.559408e-13, 1.854489e-13, 
    1.640355e-14, -6.289899e-13, -4.843972e-13, -1.113831e-13, -1.335684e-12, 
    -1.109945e-14, -4.743844e-13, 3.622797e-13, 2.173854e-13, 1.989658e-13, 
    -6.904893e-13, -2.731773e-13, -1.899349e-12, 6.003559e-13, 6.481988e-12, 
    1.274415e-13, 7.71605e-14, -5.283593e-13, 1.296826e-12, -1.047259e-13, 
    2.144951e-13, 4.64008e-12, -1.596553e-12, 1.707662e-14, -3.03866e-12, 
    3.043538e-13, 9.464651e-15, -6.609852e-13, 3.985368e-13, 1.028316e-13, 
    -2.031986e-13, 2.174233e-13, -8.100326e-13, -3.175654e-13, -1.541406e-13, 
    1.563236e-12, 1.625644e-13, 4.635459e-13, 1.597056e-13, -5.529216e-13, 
    -4.111475e-12, 1.377886e-12, 2.997366e-12, -1.690817e-11, -2.166045e-13, 
    4.32647e-13, 6.279945e-13, 4.928002e-14, -9.200141e-13, -2.019218e-14, 
    3.824441e-13, -1.326023e-13, -7.23116e-13, -1.290228e-12, -5.843243e-14, 
    -7.963075e-14, -2.837577e-12, 2.289072e-13, 1.425707e-13, -1.876554e-13, 
    -8.428064e-13, 3.763101e-14, -1.859207e-13, -1.632666e-12, -3.562067e-13, 
    -1.054934e-12, -1.024779e-12, 2.392826e-13, -6.733763e-14, -5.866002e-13, 
    5.731526e-15, 4.060641e-14, 3.222145e-13, 6.254441e-13, 1.242256e-12, 
    1.067091e-12, 8.276713e-13, 3.631262e-13, 1.688927e-13, 2.602502e-13, 
    1.982062e-12, -2.199374e-12, -2.403761e-12, 1.071712e-14, -2.05877e-13,
  5.256628e-13, 3.581857e-13, 2.868816e-13, 2.189915e-13, 2.051415e-13, 
    3.089751e-13, 1.198763e-13, -2.779443e-13, -5.657141e-13, -2.38698e-13, 
    2.345901e-13, 1.357248e-13, -5.452028e-13, 3.407552e-13, 1.375566e-13, 
    2.790518e-13, 1.856959e-13, -3.697737e-13, 2.092528e-13, 4.668765e-13, 
    5.298539e-13, 8.59951e-13, 7.950307e-13, -7.769341e-13, -7.814027e-13, 
    -1.62978e-12, 1.959266e-13, 5.639933e-14, -1.35808e-13, -9.70779e-13, 
    -7.421841e-14, 4.980738e-13, 9.121037e-13, -9.381385e-14, -1.238176e-12, 
    1.640355e-14, -6.103229e-13, 2.077651e-12, 5.781209e-13, 3.933409e-13, 
    7.258805e-13, 6.486478e-14, 6.137799e-13, 2.631688e-13, 9.878487e-13, 
    -1.909667e-12, -3.134298e-13, 1.1674e-12, 1.576222e-12, 2.11065e-11, 
    6.717474e-13, -2.696315e-12, 1.218969e-13, -9.426404e-13, -2.819196e-13, 
    -9.326706e-13, 1.580763e-12, -1.695005e-13, 3.70981e-14, -2.926812e-12, 
    -2.592371e-13, -2.803591e-13, -3.503586e-13, 2.693179e-13, 1.506739e-13, 
    6.751544e-13, -5.147549e-13, -3.302913e-13, 4.75231e-13, 5.893064e-13, 
    5.716816e-13, -3.713141e-13, 9.167112e-13, 6.413481e-13, -8.761686e-13, 
    -2.781136e-12, 1.159496e-12, -1.290287e-12, 1.143632e-12, 8.087142e-13, 
    9.257595e-13, 6.748574e-13, -1.77941e-13, -1.925793e-12, -1.289774e-12, 
    -3.644307e-14, -6.829259e-13, -5.463408e-13, 1.666054e-13, -2.95608e-12, 
    -5.074274e-13, -7.41196e-13, 2.25521e-13, 1.621631e-12, 8.842926e-13, 
    6.341708e-12, 1.169653e-12, -4.24577e-13, -1.60566e-12, 8.160528e-13, 
    -2.441158e-12, 7.872054e-13, 3.91449e-13, 4.182731e-13, 1.015854e-14, 
    -1.149081e-13, -9.917067e-14, 3.801959e-13, 1.01244e-12, 1.205452e-12, 
    1.134204e-12, 1.259742e-12, -1.125489e-13, 1.237621e-13, -5.939971e-13, 
    2.440886e-12, 1.319757e-11, -1.370819e-11, -6.409526e-13, 1.763034e-13,
  1.023764e-13, -1.083994e-13, -1.693506e-13, -1.057904e-13, -1.718486e-13, 
    -6.756679e-13, -4.701101e-13, 2.095685e-13, 5.577344e-13, 9.531403e-13, 
    -1.923323e-13, 7.190082e-14, 3.302497e-13, 1.711034e-12, -1.839501e-13, 
    7.700812e-13, 4.159645e-13, 3.930883e-13, 6.007694e-13, 4.300033e-13, 
    -1.602468e-13, 2.011294e-12, 3.564163e-12, 2.075742e-12, -3.860107e-13, 
    8.714834e-13, 1.584247e-12, 6.343398e-13, 1.242798e-12, -5.729722e-13, 
    -3.022846e-12, -8.716777e-13, -2.673181e-12, -1.982164e-13, -2.11052e-12, 
    2.595285e-13, -6.387585e-13, 2.462544e-13, 1.486603e-12, -2.018061e-12, 
    8.453932e-13, -3.382614e-12, 1.03452e-12, 7.02877e-13, -1.060527e-12, 
    -5.2338e-12, -3.805706e-13, 1.565234e-12, 3.980086e-12, 9.004283e-12, 
    1.176073e-13, -3.955933e-12, 2.120751e-12, 4.785764e-12, 5.904694e-13, 
    -6.360329e-13, -4.855422e-13, -2.001482e-13, 1.932479e-12, 1.05646e-12, 
    2.862724e-12, -3.295628e-12, -6.477457e-13, 6.514484e-13, 2.777473e-13, 
    -3.462508e-14, 5.891121e-14, -3.550424e-12, -1.532316e-12, 2.901152e-13, 
    -2.398901e-12, -2.643039e-12, 2.02395e-12, -1.64789e-12, -1.100028e-12, 
    -2.77682e-12, 1.953299e-14, -2.915446e-13, -7.435916e-12, -1.255537e-12, 
    1.473197e-12, -1.19703e-12, -5.416084e-13, -6.454143e-13, -1.236164e-12, 
    -1.064357e-12, -3.853626e-12, -8.490847e-13, -1.477364e-12, 
    -2.028516e-13, -8.868878e-13, -1.881911e-13, 2.013667e-14, -1.871559e-14, 
    1.104811e-13, -4.695952e-12, -4.894502e-13, -3.40214e-13, 5.65839e-13, 
    -4.901385e-13, -3.87633e-12, 1.885055e-12, 3.857123e-13, -7.237318e-12, 
    -5.901252e-13, -2.295247e-13, 1.229711e-13, 1.462344e-12, 1.873404e-12, 
    1.451964e-12, 4.211215e-13, 1.371583e-12, -1.097317e-13, 1.184566e-12, 
    -1.506989e-13, 1.05406e-12, 1.021281e-11, -1.857294e-12, 3.272244e-13, 
    -1.312769e-12,
  -7.132073e-13, 1.575406e-13, 1.225131e-13, 2.354783e-13, 2.161493e-12, 
    1.597833e-12, 2.59226e-12, 3.026579e-12, 5.939693e-12, 2.473466e-12, 
    3.999634e-12, 2.844669e-12, -1.303402e-13, 4.090284e-12, 9.421131e-12, 
    1.750611e-12, -1.939726e-13, 1.581013e-12, 6.902812e-13, 5.582201e-13, 
    1.238898e-12, 1.747991e-12, 2.222111e-12, 2.777722e-12, 1.050771e-12, 
    1.244688e-11, 1.130768e-11, 1.248279e-12, 3.319289e-12, 3.268164e-12, 
    2.741141e-12, 3.568257e-12, -2.526979e-12, -2.476297e-12, -6.821488e-12, 
    6.106227e-16, 2.98378e-13, 3.011688e-13, 1.929734e-12, 2.850803e-12, 
    -5.89806e-13, 5.978107e-12, 1.847272e-13, 2.12236e-12, -3.403167e-12, 
    -1.322165e-12, 1.882106e-13, -9.383466e-13, 4.51088e-12, 2.832304e-12, 
    2.775988e-12, -1.807665e-12, -7.80287e-13, 1.061828e-11, 7.974107e-13, 
    -1.884881e-13, 1.831868e-15, 3.112233e-13, 3.223921e-13, 2.958522e-12, 
    4.54381e-12, 4.899414e-13, -7.375989e-12, 1.402323e-13, -2.498668e-13, 
    1.091793e-12, -1.080069e-11, 4.692358e-13, -4.3196e-12, 1.093814e-11, 
    -5.178136e-12, -2.719769e-12, -4.048983e-13, -9.654499e-13, 
    -2.947259e-12, -2.387646e-12, -1.892445e-13, 4.199419e-13, -1.409122e-11, 
    -2.606193e-12, 2.015998e-12, 5.977899e-13, -5.424272e-13, 1.416289e-11, 
    6.010747e-13, 3.352874e-13, -1.130918e-11, 7.669421e-13, -1.267149e-12, 
    2.361972e-12, 5.635492e-13, -4.564793e-13, -1.018907e-13, 1.031453e-13, 
    3.263945e-12, -1.182953e-11, -2.037226e-12, -7.252532e-13, 2.452372e-12, 
    2.345968e-12, -2.682299e-13, 1.540667e-12, 4.042877e-13, -2.236044e-11, 
    -8.724133e-13, -3.591571e-14, 3.926859e-13, 1.343203e-12, 9.599543e-13, 
    9.610646e-13, 9.289791e-13, 2.551959e-12, 2.507106e-12, 1.096012e-12, 
    -2.431944e-12, 3.695155e-13, 1.142163e-12, -3.150891e-12, 2.91444e-13, 
    2.538636e-12,
  -1.553757e-13, 3.278544e-12, 3.394229e-12, 6.999512e-12, 1.099476e-11, 
    8.626488e-12, 1.056161e-11, 6.265766e-12, -3.943179e-12, 2.192246e-12, 
    5.170642e-12, 2.043976e-12, 3.67939e-12, -3.230305e-12, 2.462919e-12, 
    3.387901e-12, 2.004757e-12, -4.490713e-12, -9.834356e-13, 3.890832e-12, 
    3.242295e-12, 1.387057e-12, 3.897993e-13, -3.911871e-13, 1.08204e-11, 
    2.135697e-11, 2.470796e-11, 9.717449e-12, 3.70548e-12, -8.512635e-13, 
    8.973378e-13, 3.169964e-12, 1.932898e-12, -6.420531e-12, -2.260192e-12, 
    -6.086742e-12, -1.411149e-12, 5.722922e-13, 3.036071e-12, 3.612777e-13, 
    1.674272e-12, 6.64141e-12, 2.261066e-12, 1.799534e-12, -4.173994e-12, 
    7.958079e-12, 1.81774e-12, 2.960132e-13, 4.958567e-12, -9.051732e-12, 
    7.311325e-12, 2.626233e-13, 5.458245e-13, 4.264589e-13, 3.028577e-13, 
    -2.571832e-13, -4.512835e-12, 1.121719e-12, -3.689687e-12, 3.148849e-12, 
    -5.534462e-13, 1.351702e-11, -4.898359e-12, 4.319212e-12, 2.178291e-12, 
    -9.471496e-11, -3.810946e-11, -7.351675e-12, 6.702694e-12, -6.517342e-12, 
    -1.695977e-12, -1.548373e-12, -4.26853e-12, -4.286016e-13, -8.688266e-12, 
    -1.150524e-12, -1.3365e-13, 5.501155e-13, -1.072864e-11, 3.054668e-12, 
    3.934741e-12, -1.94959e-11, 1.878914e-12, 2.485179e-11, 6.054601e-13, 
    -1.280198e-12, -1.08849e-11, 3.099188e-13, 1.929716e-12, -6.586953e-13, 
    1.697753e-12, 9.063971e-13, -3.319567e-14, 1.691935e-12, 7.519763e-12, 
    -6.513129e-12, -4.643197e-12, -1.772582e-12, 2.143785e-12, 3.457845e-12, 
    2.382372e-12, 2.731131e-12, -8.655923e-14, -4.721482e-11, 4.28102e-13, 
    1.021017e-12, -1.295353e-12, 1.551759e-12, 6.413758e-13, -2.399192e-13, 
    3.07393e-12, 7.01772e-13, -1.653844e-12, -4.821032e-12, 4.010681e-13, 
    4.80227e-14, -4.665018e-14, -4.711939e-12, -9.528489e-14, 1.359624e-11,
  -3.928385e-13, 1.297552e-11, 6.912818e-12, 5.595371e-12, 1.387571e-12, 
    2.643732e-12, -1.166643e-11, 4.51887e-11, 6.432362e-11, 2.906304e-11, 
    1.877901e-12, 4.316131e-13, -6.717266e-13, -5.696041e-12, -9.445486e-12, 
    3.825343e-12, 1.336828e-12, -6.471754e-12, 4.281644e-13, 3.264847e-12, 
    1.939143e-13, -2.798636e-12, -3.131093e-12, -1.425808e-11, 2.468206e-12, 
    -6.619864e-11, -4.093763e-11, 1.034008e-11, -2.724085e-12, -3.395437e-12, 
    4.639414e-12, -1.351556e-11, -4.455422e-12, -4.959574e-12, 1.254281e-11, 
    5.174264e-12, -8.111742e-12, 3.010092e-13, 9.052883e-12, -3.179376e-12, 
    1.097613e-11, -4.11754e-14, -1.897649e-13, -4.652433e-13, 2.253489e-12, 
    6.580528e-12, 4.059156e-12, 2.592385e-12, 8.136017e-12, -8.739457e-12, 
    1.635872e-12, -1.983275e-13, 8.265888e-14, -6.312589e-13, 4.409015e-13, 
    1.406791e-13, -3.157016e-12, 2.660508e-12, -1.348602e-12, 1.955334e-11, 
    -1.152249e-11, 3.869252e-12, -3.583842e-12, -8.33908e-13, -3.500575e-12, 
    -3.749927e-11, 8.840845e-13, -6.254858e-13, -8.327089e-13, 3.59396e-11, 
    1.488823e-12, -5.633265e-11, 4.598669e-12, -1.982441e-11, -6.730991e-12, 
    -2.096517e-13, -3.504419e-13, 4.377054e-14, 4.388979e-12, 8.661252e-12, 
    9.801174e-12, -5.955127e-11, 2.422132e-12, 1.060514e-11, -6.824749e-12, 
    -3.956876e-12, -2.447806e-12, -6.265918e-12, 1.322696e-12, -1.289011e-12, 
    5.319481e-12, -9.363119e-12, -3.264888e-13, 2.341929e-12, 2.604167e-13, 
    -4.72383e-12, 3.614234e-12, -1.827136e-12, -2.170361e-12, 3.989156e-12, 
    -7.307308e-12, 2.16337e-12, -3.705473e-13, -3.4243e-11, 7.154971e-13, 
    1.055281e-12, -3.400044e-12, -9.982432e-13, -6.686734e-13, 2.212744e-12, 
    -1.97313e-12, -4.159381e-12, -5.617493e-12, 1.586412e-12, 2.355408e-12, 
    -3.851336e-13, 4.377748e-14, -3.819873e-12, 1.749399e-13, 4.093573e-12,
  -2.785328e-12, 1.935119e-12, 2.90834e-12, 7.224221e-12, 3.810174e-12, 
    1.911693e-12, 1.004314e-10, 3.572859e-11, -5.892975e-11, -5.56164e-11, 
    -3.810952e-12, -3.047007e-12, -9.836687e-12, 8.414269e-12, -2.061407e-12, 
    -9.178879e-13, -1.38668e-12, -5.128231e-12, -2.389616e-13, 5.605738e-12, 
    1.266609e-11, 2.454331e-11, 2.682771e-11, -2.489298e-11, 4.172107e-12, 
    3.477779e-11, 4.281131e-12, 1.765615e-11, -3.487211e-13, -3.702011e-11, 
    1.60843e-11, 6.204648e-12, 2.607858e-12, -8.163803e-12, 5.857981e-12, 
    2.025391e-11, -2.976769e-12, 7.85344e-14, 1.99743e-11, -2.030664e-12, 
    2.031464e-12, -1.23257e-12, 5.625223e-12, -1.28803e-12, 4.931167e-12, 
    9.197088e-12, 4.005019e-12, 5.300677e-12, 9.692314e-12, -1.789079e-12, 
    -6.68389e-13, -2.154943e-13, -5.931922e-13, 7.795986e-14, -5.262832e-13, 
    4.962142e-13, 3.645084e-12, 1.984324e-12, -3.088707e-12, 1.831112e-11, 
    -2.752126e-11, 1.267431e-12, 1.009637e-12, -4.774681e-12, -7.779677e-12, 
    -1.388473e-11, 6.809109e-12, 7.051476e-11, -6.534689e-11, 4.328493e-11, 
    -3.008543e-11, 7.592371e-12, 1.351191e-11, -1.926626e-12, 6.63819e-12, 
    -2.368661e-12, -7.793211e-13, 3.272688e-12, 1.159791e-11, 8.295031e-13, 
    7.801371e-12, -8.680759e-12, 5.598577e-13, 4.248296e-11, -5.626832e-12, 
    8.286705e-13, 6.539935e-12, -8.15864e-12, -3.001219e-13, -8.74828e-13, 
    4.581391e-12, -1.160232e-11, -9.256901e-13, 5.397266e-12, 7.031598e-13, 
    -1.967554e-12, 2.430078e-12, 8.135881e-12, -2.824019e-12, 2.427658e-12, 
    -1.260131e-11, 5.675977e-12, -3.234982e-13, -2.489176e-12, -8.086865e-13, 
    3.054945e-12, 2.392531e-12, -3.146317e-12, -4.323264e-12, 3.224365e-12, 
    -1.215267e-11, -9.373058e-12, 4.465484e-12, 2.094208e-11, -3.447131e-12, 
    -1.370681e-13, 7.935319e-14, -2.184542e-12, 2.547046e-12, 3.163247e-12,
  -8.386847e-12, 1.181499e-12, 1.169498e-11, 2.38638e-11, 5.224332e-11, 
    1.353792e-10, 6.262479e-11, -7.73992e-12, -9.569523e-11, -2.959655e-11, 
    -1.997502e-11, -1.059752e-11, -5.970002e-12, 1.970923e-11, 1.565326e-11, 
    -2.21323e-12, -3.673983e-12, -5.404954e-12, -1.12392e-12, 8.94218e-12, 
    7.661871e-12, -1.175382e-11, 2.870271e-11, -9.220513e-12, 5.716616e-11, 
    -2.017941e-12, 1.52246e-11, -3.06678e-11, -1.117295e-11, -1.787914e-11, 
    8.961054e-12, -2.003986e-11, 2.149214e-11, -1.163203e-11, -1.078793e-11, 
    -7.448642e-11, -3.811396e-13, -3.390344e-14, 6.306622e-12, 3.540168e-13, 
    4.966161e-12, 1.493816e-11, 4.704404e-12, -1.877866e-12, 1.615563e-11, 
    -7.778667e-12, 4.553968e-12, 6.286638e-12, 5.889267e-12, 1.950939e-13, 
    1.990907e-13, -2.038791e-11, -4.083733e-13, 1.36251e-12, 3.159667e-13, 
    3.251288e-13, 6.148304e-12, 8.150147e-13, -1.296452e-12, 1.66825e-11, 
    -2.805656e-11, 3.043343e-12, 8.484324e-13, -4.966294e-12, -6.016876e-12, 
    -7.957845e-11, 1.572076e-13, 7.829826e-11, 3.296441e-11, 3.43533e-11, 
    -3.283007e-11, -1.250011e-11, 5.359357e-11, 9.291456e-13, 4.622936e-12, 
    -3.327671e-12, -8.725937e-13, 6.836642e-12, 6.211559e-13, 7.127743e-12, 
    3.560263e-12, 8.797904e-11, 2.303713e-14, 5.524869e-11, 1.39827e-11, 
    4.063994e-11, -2.764367e-11, -2.137401e-12, -1.021081e-12, -6.178391e-13, 
    2.167266e-12, -1.427585e-11, -1.760814e-12, 7.129553e-12, -2.807166e-11, 
    -6.355561e-12, 1.01148e-12, 2.185252e-11, -1.625711e-11, -1.639289e-12, 
    -2.155343e-11, 5.161913e-13, 8.484879e-14, 9.964217e-12, -1.971345e-11, 
    1.088463e-12, -2.319145e-12, 2.010503e-12, 1.205414e-11, 3.3058e-12, 
    -1.400868e-11, -7.213674e-12, 5.2367e-12, 2.45266e-11, -5.583534e-12, 
    -2.107203e-14, 2.812611e-13, -7.817184e-13, 1.051936e-11, 5.575651e-12,
  -9.205081e-12, -4.825917e-12, 4.483747e-11, 1.243439e-10, 1.091345e-10, 
    6.431988e-11, 7.633671e-12, -3.765876e-11, -1.248379e-11, 1.181886e-10, 
    -1.549494e-11, -6.631451e-11, 8.371748e-12, -1.085398e-11, 2.917933e-11, 
    -1.398615e-12, -4.735123e-12, -3.038791e-12, -2.978451e-12, -1.00675e-12, 
    -8.86935e-12, -2.202682e-12, 4.669065e-11, -1.972511e-11, 4.329026e-11, 
    1.056788e-10, 2.688694e-11, -9.523426e-11, -4.885647e-12, 1.613842e-11, 
    3.256284e-11, -4.900969e-12, 1.874145e-11, -1.18705e-12, 8.116396e-12, 
    -2.33783e-10, -2.871014e-12, -9.517387e-14, -6.45084e-12, 5.14544e-13, 
    -2.751577e-13, 2.484835e-11, -6.0843e-12, -2.497239e-13, -2.042588e-12, 
    -3.108624e-11, 3.939626e-12, 4.346301e-12, -6.921574e-13, -9.686696e-15, 
    7.908896e-12, -5.6257e-11, 4.710899e-13, 9.217072e-13, 1.57343e-12, 
    -5.322409e-13, -1.163492e-11, 3.690825e-13, 3.386469e-12, -2.034262e-11, 
    -2.472911e-11, 1.526557e-12, -1.565414e-12, -4.08189e-12, -3.577982e-12, 
    1.025275e-10, -3.069034e-11, 1.806746e-10, -4.24567e-11, -1.637357e-12, 
    -3.141665e-11, 1.153522e-12, 5.643308e-11, -1.02891e-11, -1.723022e-12, 
    -7.66498e-13, -4.995726e-13, -3.838374e-12, -7.486456e-13, 1.613798e-11, 
    3.713696e-13, 9.766653e-11, 2.308154e-13, 5.384004e-11, -8.334555e-11, 
    4.769518e-11, 4.148171e-11, 1.059042e-11, -1.039134e-13, -1.065925e-12, 
    -2.715383e-11, -1.855027e-11, -1.703415e-12, -1.660438e-11, 
    -6.657275e-11, -7.925771e-12, -8.988588e-12, 1.033174e-12, -1.604095e-11, 
    -4.166223e-12, -8.133494e-12, -1.303679e-11, 1.205869e-12, 7.945589e-13, 
    -2.98892e-11, -6.616929e-13, 8.499867e-13, 3.395018e-11, 2.716338e-11, 
    3.804734e-12, -8.638201e-12, -3.86069e-12, -1.467049e-12, 8.168355e-12, 
    4.442224e-12, -6.386003e-14, 2.312595e-13, 1.094402e-12, 9.634002e-12, 
    -8.889334e-12,
  -6.479572e-11, 2.568812e-11, 1.249594e-10, 1.321658e-10, 1.278488e-11, 
    -1.42053e-11, -3.944955e-11, 1.130254e-10, 3.289893e-10, 1.913689e-10, 
    -2.475482e-10, -8.07161e-11, 1.530183e-10, -4.916401e-11, -3.13376e-11, 
    -2.007727e-13, -4.602918e-12, -3.192224e-12, -8.541667e-12, -3.98015e-12, 
    1.444622e-12, 9.333201e-12, 3.216005e-11, -5.972112e-12, -7.586376e-12, 
    2.592024e-10, -1.810463e-11, -4.581313e-11, 2.995604e-12, 3.251199e-11, 
    4.344769e-11, 8.220979e-12, 1.003042e-10, 3.753886e-11, 6.313305e-11, 
    1.189193e-10, -1.518297e-12, -1.731393e-13, 7.617307e-11, 2.998046e-13, 
    -9.895595e-12, 2.236988e-11, -3.764933e-12, 2.274313e-12, -4.900058e-11, 
    1.227218e-11, 3.671508e-12, 2.082945e-12, -2.315525e-12, 2.553513e-13, 
    2.225256e-11, -5.797007e-11, -8.248735e-13, 1.911626e-12, 7.412404e-13, 
    -3.604894e-13, -2.043921e-11, -6.623591e-13, 2.642353e-12, -6.375844e-12, 
    -3.003153e-11, 1.333755e-11, -1.654188e-11, -4.553691e-12, -2.768585e-12, 
    5.075349e-10, -1.063714e-10, 4.628369e-10, -2.676415e-11, -6.993739e-12, 
    4.706235e-12, -5.07594e-12, 9.84679e-11, -4.764078e-11, 1.039457e-12, 
    9.503509e-14, -1.085243e-13, -2.549572e-12, -2.647471e-12, 2.71394e-11, 
    -3.454459e-12, 4.615168e-11, 1.026623e-12, 7.656098e-11, -5.021739e-11, 
    7.242784e-11, 9.62288e-11, 2.908584e-11, 4.359534e-13, -3.069767e-13, 
    -4.211764e-11, -9.078516e-12, -5.061507e-13, -5.150867e-11, 
    -1.073612e-10, -1.13862e-11, -7.914825e-12, -7.181877e-11, -1.915246e-11, 
    -3.157341e-12, 1.202372e-11, -9.385145e-12, 1.965872e-12, -5.841161e-14, 
    -1.66327e-11, 2.087153e-11, 3.953793e-11, 3.262857e-11, 2.302381e-12, 
    6.042722e-12, -2.438272e-12, -2.541301e-12, -1.713163e-11, -8.703926e-12, 
    2.66025e-11, -4.070078e-14, -8.337775e-14, 1.298843e-12, 4.034342e-12, 
    -9.201084e-12,
  -9.936163e-11, 6.845347e-11, 1.24069e-10, 2.613487e-11, -5.735123e-11, 
    -5.117662e-11, 2.130274e-11, 2.765852e-10, 3.95699e-11, -2.915057e-10, 
    -4.484346e-11, -1.262819e-10, 1.379112e-10, -9.70648e-11, -5.797607e-11, 
    -8.228973e-14, -4.819966e-12, -2.922773e-12, -1.072964e-11, 8.565815e-12, 
    1.823852e-11, 3.097189e-11, -9.419798e-12, -1.761635e-11, -9.186207e-12, 
    3.101766e-10, 1.804563e-10, -1.834377e-11, 4.943379e-12, -6.010081e-12, 
    7.318968e-11, 1.008742e-10, -7.707235e-11, 4.43785e-11, 9.355294e-11, 
    3.577869e-10, 1.63829e-12, -1.636469e-13, 1.510607e-10, -1.132872e-13, 
    -3.551688e-11, 2.173439e-11, 8.899548e-12, -9.294995e-13, -9.753598e-11, 
    3.559086e-11, 4.343859e-12, 8.951728e-13, -6.834666e-12, 1.514955e-12, 
    3.390455e-11, -5.330913e-11, -2.966072e-12, 1.603295e-12, 1.776024e-13, 
    3.439471e-13, 1.730667e-10, -4.356959e-13, -9.880719e-12, 1.97114e-11, 
    -5.196665e-11, 3.571521e-11, -4.742984e-11, -4.552581e-12, -3.944711e-12, 
    3.184983e-10, 1.147489e-10, 5.018441e-10, -2.864486e-11, 1.812039e-11, 
    -8.344592e-11, 5.248313e-11, -1.536793e-11, -4.893397e-11, 1.440905e-11, 
    4.500844e-13, -3.441691e-15, 9.122703e-12, -4.700318e-12, 4.885181e-11, 
    -5.31819e-12, 3.038038e-11, 1.585398e-12, -5.410361e-11, 9.696621e-11, 
    1.860043e-10, 1.355012e-10, 4.582756e-11, 1.46913e-12, 3.936185e-12, 
    -3.600653e-11, -4.164624e-12, 5.571099e-13, -3.289915e-11, -1.392075e-10, 
    -1.157643e-11, 5.406476e-12, -3.267542e-11, -4.783929e-11, -2.637135e-12, 
    1.954681e-11, 1.789235e-12, 2.343514e-12, 1.916522e-13, -2.017386e-11, 
    -2.458767e-11, -5.633605e-11, -1.587819e-11, -9.311441e-12, 1.292899e-11, 
    -3.254064e-12, -2.723821e-12, -3.451306e-11, -3.581357e-12, 4.322964e-11, 
    6.639134e-14, 5.040413e-14, 1.542239e-13, 2.253864e-12, 6.034129e-11,
  -8.586376e-11, 7.02034e-11, 6.650946e-11, -6.639045e-11, -4.3066e-11, 
    8.072121e-11, 1.700249e-10, 9.050805e-11, 1.551044e-10, -3.224807e-10, 
    1.192113e-11, -1.222897e-10, -5.311396e-11, -1.369003e-10, -1.091642e-10, 
    5.870859e-14, -5.065815e-12, -3.9031e-12, 8.888446e-13, 3.612932e-11, 
    2.016698e-11, 3.697576e-11, -7.476952e-11, -4.174741e-10, -6.388223e-11, 
    3.015739e-10, 3.797931e-10, -3.864375e-11, -8.330403e-11, -1.901066e-10, 
    -7.092193e-11, 7.624923e-11, 8.355183e-11, 3.06386e-11, 1.709184e-10, 
    4.594733e-10, 5.306067e-12, -1.163514e-13, 1.245057e-10, -1.485034e-13, 
    -8.869421e-11, 1.145573e-11, 1.948552e-11, -4.617737e-12, -3.218199e-10, 
    -5.078959e-11, 8.817835e-12, 1.450839e-12, -1.433644e-11, 1.854128e-12, 
    3.692835e-11, -8.768275e-11, -2.16005e-12, -6.596323e-12, 3.306244e-13, 
    -2.362555e-13, 1.053557e-11, 1.011724e-12, -3.69373e-11, 3.533385e-11, 
    -8.276491e-11, 5.843059e-11, -5.132783e-11, -4.548717e-12, -5.290168e-12, 
    1.474074e-10, 2.692149e-10, 5.120526e-10, -5.320011e-11, 2.349498e-11, 
    -1.660085e-10, 8.315748e-11, 2.330625e-10, -6.794476e-11, 2.051603e-11, 
    -8.881784e-15, 5.928591e-14, -1.131006e-11, -3.925127e-12, 5.193534e-11, 
    -3.376854e-12, 1.791112e-11, 2.083667e-12, -1.431637e-10, 1.775167e-10, 
    3.364589e-10, -7.713385e-11, 5.955414e-11, 5.342699e-12, 1.294787e-11, 
    -3.09246e-11, 5.510436e-12, 5.719869e-13, 5.033396e-12, -1.342633e-10, 
    -3.559819e-12, 3.021903e-11, 2.84599e-11, -6.194867e-11, -4.670042e-12, 
    2.262102e-11, 2.485678e-11, 1.729894e-12, 1.472933e-12, -2.800249e-11, 
    -1.059162e-10, -1.805232e-10, -9.553602e-11, -2.673417e-12, 2.743406e-11, 
    -3.852918e-12, 2.298606e-12, -4.037659e-11, 1.403855e-11, 4.546497e-11, 
    6.030732e-14, 9.848788e-13, -3.764766e-13, 1.72351e-12, 1.551292e-10,
  -7.709211e-11, 7.099121e-11, 1.996625e-12, -6.379874e-11, 9.745271e-11, 
    1.974847e-10, 3.69802e-11, -1.698819e-10, 3.462475e-10, -3.968923e-10, 
    -3.88205e-11, -2.01239e-10, -1.834843e-10, -1.828377e-10, -1.962341e-10, 
    -4.923173e-13, -2.574296e-12, -6.75815e-12, 1.277611e-11, 5.699885e-11, 
    2.035794e-11, 5.300382e-11, -6.92042e-11, -8.751977e-10, -1.174438e-10, 
    7.652723e-11, 4.034257e-10, -6.304735e-11, -2.416876e-10, -2.215756e-10, 
    -5.471081e-10, 2.412017e-10, 6.807976e-11, 2.50572e-10, 2.608491e-10, 
    -2.547624e-10, 1.001199e-11, -1.109113e-13, 3.494849e-10, 2.657696e-12, 
    -2.502315e-10, -1.182165e-12, 1.930123e-11, -6.51354e-12, -3.433884e-10, 
    -3.579803e-11, 1.57141e-11, 5.191847e-12, -2.900666e-11, -9.677259e-13, 
    3.15995e-11, -1.993152e-10, -4.68976e-12, -1.87832e-11, 6.445289e-13, 
    -7.345236e-13, -3.664837e-10, 2.92788e-12, -7.427632e-11, -4.352407e-11, 
    -1.102158e-10, 5.923972e-11, -4.136247e-12, -7.293721e-12, -5.930367e-12, 
    1.796341e-11, 2.117684e-11, 2.116618e-11, -2.467875e-10, -1.265477e-11, 
    -1.89055e-10, 9.711076e-11, 1.05107e-10, -6.992718e-11, 1.924541e-11, 
    -1.166178e-12, 2.317035e-13, -5.053336e-11, 2.358735e-12, 4.241585e-11, 
    7.838175e-13, -1.105471e-11, 9.046097e-13, -2.910827e-10, -1.567111e-10, 
    6.922347e-10, -3.306102e-10, 6.985701e-11, 1.235106e-11, 3.461986e-11, 
    -4.594725e-11, 6.816432e-11, 1.207034e-12, 1.386917e-11, -7.228884e-11, 
    3.956302e-12, 6.029257e-11, 1.814948e-10, -4.828937e-11, -5.938184e-12, 
    1.660894e-13, 7.707879e-11, 1.449396e-13, 2.595868e-12, -8.622969e-11, 
    -9.582202e-11, -1.690168e-10, -8.397105e-11, -1.324718e-11, 3.560796e-11, 
    2.249756e-12, 7.084111e-12, -4.008083e-11, 2.031886e-11, 2.757528e-11, 
    7.727152e-14, 2.424616e-12, 1.151856e-14, 6.368239e-13, 1.924683e-10,
  -7.739764e-11, 9.306156e-11, -3.031531e-11, 3.464073e-11, 1.808331e-10, 
    7.297452e-11, -9.924861e-11, -4.284164e-10, 1.097327e-10, -7.627055e-10, 
    -3.606981e-10, -4.602345e-10, -3.415952e-10, -2.460148e-10, 
    -2.267697e-10, -1.409539e-12, 3.49889e-12, -6.820322e-12, 1.738498e-11, 
    5.509904e-11, 1.795009e-11, 8.819789e-11, 9.018564e-11, -1.250939e-09, 
    -7.426415e-11, -1.015117e-10, 2.578968e-10, -8.190959e-11, -6.401155e-10, 
    5.03082e-11, -4.499618e-10, 2.12145e-10, -4.806644e-11, 1.009576e-09, 
    1.615899e-10, -2.444729e-10, 9.910473e-12, -1.918465e-13, 4.841496e-10, 
    1.320952e-11, -4.056286e-10, -5.163514e-11, 6.859846e-12, -6.736139e-12, 
    -4.965557e-10, -1.621139e-10, 1.931877e-11, 1.631406e-11, -5.389396e-11, 
    -5.876521e-12, 2.295675e-11, -2.591012e-10, -2.420677e-11, -1.540457e-11, 
    5.577316e-13, -1.196376e-12, -3.90683e-10, 3.975131e-12, -1.168058e-10, 
    -1.834346e-10, -1.37149e-10, 2.818723e-11, 7.735856e-11, -8.368417e-12, 
    -2.99849e-13, -1.474305e-10, -4.032561e-10, -1.880629e-09, -4.278569e-10, 
    -9.547918e-11, -3.936336e-10, 8.583179e-11, -3.744649e-10, -3.156941e-11, 
    2.077041e-11, -6.387779e-12, 4.192202e-13, -7.426681e-11, 1.478897e-11, 
    4.370726e-11, 6.211032e-12, -1.438529e-11, -2.61835e-12, -3.894609e-10, 
    -4.990266e-10, 5.005703e-10, -5.688392e-10, 6.933831e-11, 2.404876e-11, 
    8.642775e-11, -1.51898e-10, -3.860272e-11, 3.887557e-12, -6.123635e-12, 
    -7.446666e-11, 1.654907e-11, 8.559766e-11, 4.319194e-10, -1.658229e-11, 
    7.648993e-13, -1.087539e-10, 2.40725e-10, -1.247003e-12, 3.620548e-12, 
    -2.473008e-10, -1.600995e-10, -1.482778e-10, 1.888445e-10, 7.328183e-11, 
    2.996181e-11, 9.942269e-12, 8.604673e-12, -3.440093e-11, 1.431211e-11, 
    -2.167155e-12, 3.078426e-13, 3.482326e-12, 1.401546e-12, -2.514766e-12, 
    1.845155e-10,
  -6.984635e-11, 1.75568e-10, 1.017266e-10, 1.389893e-10, 2.046647e-10, 
    3.574741e-11, -9.655388e-11, -5.122427e-10, -1.155897e-09, -1.498988e-09, 
    -3.396483e-10, -4.919869e-10, -2.000746e-10, -3.042189e-10, 
    -1.059686e-10, -1.215028e-12, 1.373319e-11, 2.315481e-12, 2.454059e-11, 
    4.08491e-11, 1.61986e-11, 1.063487e-10, 1.824212e-10, -1.233049e-09, 
    -1.421778e-10, -1.477911e-10, 1.73543e-10, 3.272067e-10, -8.365788e-10, 
    4.006591e-10, -5.501963e-10, -2.413181e-10, -7.131025e-10, 2.406614e-09, 
    1.986713e-10, 3.904663e-10, 2.838441e-12, 4.856116e-13, 1.200604e-10, 
    3.997425e-11, -4.468994e-10, -1.526992e-10, -7.380763e-12, -9.241941e-12, 
    -4.218172e-10, -7.589893e-10, 2.099565e-11, 4.031309e-11, -9.015935e-11, 
    -1.137401e-11, 2.374767e-12, -1.145075e-10, -7.022685e-11, -1.527312e-12, 
    1.386891e-13, -1.817213e-12, -7.493561e-10, 1.836043e-12, -2.116831e-10, 
    1.109308e-10, -1.656879e-10, -2.997069e-11, 2.604796e-10, -1.066418e-11, 
    6.743051e-13, -2.030607e-10, 2.381366e-10, -4.99417e-09, -2.683009e-10, 
    -2.865477e-10, -9.812418e-10, -1.087592e-10, -5.468319e-10, 
    -7.905321e-11, 3.311165e-11, -1.390354e-11, 3.63265e-13, -5.981482e-11, 
    3.5888e-11, 9.708856e-11, 3.040235e-12, -4.35394e-12, -6.975753e-12, 
    -6.733583e-10, -3.444711e-11, 1.61803e-10, -7.646985e-10, 5.094414e-11, 
    4.813339e-11, 2.091411e-10, -3.026877e-10, -3.028283e-10, 9.242385e-12, 
    -1.208674e-10, -1.368328e-10, 2.323049e-11, 9.007301e-11, 5.033112e-10, 
    9.602985e-12, 7.598189e-12, -1.610587e-10, 4.693838e-10, -1.084022e-12, 
    9.123258e-12, -5.17387e-10, -4.304468e-10, -3.957314e-10, 7.621406e-10, 
    5.762146e-10, 3.017675e-11, 1.693934e-11, 2.384226e-11, -6.470735e-11, 
    -2.273914e-11, -3.194423e-11, 1.098499e-12, 4.838352e-12, 3.454848e-12, 
    -6.450285e-12, 1.534914e-10,
  -1.294289e-10, 3.337952e-10, 4.299636e-10, 3.059064e-10, 3.235705e-10, 
    2.293028e-10, -1.402114e-10, -6.528467e-11, -1.86451e-09, -2.163386e-09, 
    2.004263e-10, 4.68809e-10, -9.706724e-11, -3.232827e-10, -2.485692e-10, 
    -7.460343e-12, 2.392007e-11, 2.593126e-11, 3.578826e-11, 3.211653e-11, 
    2.381384e-11, 9.585222e-11, 1.122338e-10, 2.633804e-10, -3.782965e-10, 
    -1.171365e-10, 3.212506e-10, 5.455512e-10, -9.219683e-10, 2.075314e-09, 
    4.645884e-10, -7.707506e-10, -1.546503e-09, 4.1356e-09, 1.572573e-10, 
    6.984635e-12, -2.646381e-11, 3.500311e-12, -2.617782e-10, 8.171028e-11, 
    -7.771845e-11, -2.258638e-10, 8.828493e-13, -1.997924e-11, -5.463257e-10, 
    -1.609596e-09, 4.649614e-11, 8.911893e-11, -9.92209e-11, -2.059175e-11, 
    -4.320988e-13, 4.85656e-12, -1.451138e-10, 1.969696e-11, 5.230039e-12, 
    -2.000178e-12, -8.014851e-10, -5.600497e-12, -4.802835e-10, 1.056133e-10, 
    -2.166658e-10, -8.375878e-11, 2.302443e-10, -1.587637e-11, -1.209131e-11, 
    -3.394263e-11, 6.332783e-10, -4.060304e-09, -8.337508e-11, -5.764029e-10, 
    -1.489319e-09, 2.352643e-10, -4.809984e-10, -2.644107e-10, 4.062173e-11, 
    -1.907807e-11, -7.700507e-13, -2.54472e-11, 5.767067e-11, 1.284981e-10, 
    -2.332712e-11, 1.490265e-10, -1.44631e-11, -7.557439e-10, 8.703012e-10, 
    -5.723777e-10, -6.672067e-10, 2.495781e-11, 1.201619e-10, 4.987228e-10, 
    -6.22375e-10, -3.20319e-10, 1.378542e-11, -2.851436e-10, -1.740013e-10, 
    -6.647482e-12, 7.897043e-11, 3.624301e-10, 4.158807e-11, 1.62224e-11, 
    3.645795e-11, 5.870981e-10, 6.119549e-12, 2.900014e-11, -7.114345e-10, 
    -7.80247e-10, -6.836025e-10, 1.13614e-09, 1.616716e-09, 1.141167e-10, 
    1.905676e-11, 4.604672e-11, -8.940759e-11, -7.814549e-11, -6.842527e-11, 
    3.64615e-12, 7.243983e-12, 4.67737e-12, -7.229994e-12, 1.041975e-10,
  -1.431211e-10, -1.371703e-11, 5.555982e-10, 4.967013e-10, 4.694165e-10, 
    3.974741e-10, 8.848033e-11, 3.254605e-10, -1.461668e-09, -1.897792e-09, 
    1.873026e-10, -2.062102e-10, 7.072565e-10, -3.248637e-10, -1.862581e-10, 
    -7.984795e-11, -3.550582e-12, 6.399503e-11, 4.763923e-11, 3.611333e-11, 
    5.423928e-11, 5.105605e-11, 7.840484e-11, 1.669232e-09, -3.276703e-10, 
    3.318839e-10, 1.678124e-10, 2.850804e-10, -7.158043e-10, 3.438348e-09, 
    3.213749e-10, -1.179867e-09, -1.666148e-09, 5.876498e-09, 3.640466e-11, 
    -1.582624e-09, -7.480167e-11, 7.96696e-12, -1.486672e-09, 1.255529e-10, 
    -1.448818e-10, -1.831388e-10, 6.185807e-11, -6.155654e-11, -6.318466e-10, 
    -1.333422e-09, 1.206146e-10, 2.52367e-10, -1.033577e-10, -3.721912e-11, 
    1.414984e-10, 1.812772e-10, -1.643528e-10, 1.062141e-10, 2.878604e-11, 
    -1.03384e-12, 3.958789e-11, -1.786802e-11, -1.116846e-09, -3.004033e-10, 
    -2.755023e-10, -1.35902e-10, -7.589662e-11, -1.250626e-11, -2.289013e-11, 
    2.789982e-10, 1.436856e-09, -3.786194e-09, -2.32372e-09, -8.620624e-10, 
    -1.130172e-09, 1.028983e-09, -3.100986e-10, -7.865246e-10, 6.365397e-11, 
    -1.144329e-11, -3.311129e-12, 1.889155e-11, 6.525767e-11, -2.80675e-10, 
    -5.680079e-11, 5.810832e-10, -2.935963e-11, -5.489973e-10, -7.386447e-11, 
    -1.512976e-09, -1.880842e-10, 6.348699e-12, 3.949676e-10, 9.405561e-10, 
    -1.315019e-09, -3.124988e-10, 1.363176e-11, -4.159375e-10, -1.748823e-10, 
    -7.237375e-11, 1.0509e-10, 2.082423e-10, 2.29825e-11, 4.044622e-11, 
    1.127276e-11, 5.997296e-10, 1.903011e-11, 6.590994e-11, -6.984742e-10, 
    -9.052705e-10, -7.2394e-10, 6.319674e-10, 2.304301e-09, 4.573941e-10, 
    -2.34941e-11, -1.817924e-11, -5.286793e-11, -1.155662e-10, -1.177263e-10, 
    8.505907e-12, 1.159695e-11, 3.274048e-12, -8.510526e-12, 3.683809e-11,
  -1.222489e-10, -6.492016e-10, 8.264536e-10, 1.325766e-09, 2.484697e-10, 
    4.630536e-10, 7.082477e-10, 8.723333e-11, 1.363887e-10, -1.043041e-09, 
    -6.016236e-10, 8.434853e-11, -1.115531e-09, -3.411529e-10, -1.736638e-10, 
    -2.928033e-10, -2.430283e-10, 9.702461e-11, 2.755307e-11, 7.89484e-11, 
    1.207852e-10, 5.179857e-12, 1.191509e-10, 2.362533e-09, -2.864148e-09, 
    2.047251e-09, -9.057359e-10, -9.685053e-10, -8.593943e-10, 3.092772e-09, 
    -1.701089e-09, -2.034049e-09, -1.936264e-09, 7.841187e-09, 9.722356e-11, 
    3.378837e-09, -7.201067e-11, 1.234746e-11, -1.708223e-09, 1.559442e-10, 
    -1.405894e-10, -9.682566e-11, 9.089973e-11, -2.441367e-10, -5.422081e-10, 
    -2.806431e-10, 2.153939e-10, 6.627801e-10, -1.877069e-10, 1.615685e-11, 
    5.684129e-10, -2.05894e-10, -5.832419e-11, 2.289667e-10, 5.014122e-11, 
    1.058709e-12, 1.30057e-09, -3.14941e-11, -2.127058e-09, -5.946177e-10, 
    -3.146923e-10, -2.050129e-10, -1.78467e-10, 9.050894e-12, -2.394955e-11, 
    2.36701e-09, 1.393374e-11, 2.780993e-10, -1.333298e-09, -8.409913e-10, 
    6.362555e-10, 1.936307e-09, -2.273026e-11, -1.132342e-09, 5.944685e-11, 
    9.883649e-12, -4.714451e-12, 6.418333e-11, 3.626397e-11, -4.127898e-10, 
    -2.196998e-11, 1.072418e-09, -5.409362e-11, 8.004193e-10, -9.498322e-10, 
    -3.96021e-10, 1.165795e-09, -1.58451e-12, 1.032729e-09, 1.177064e-09, 
    -2.427406e-09, -3.232756e-10, 9.64917e-12, -1.785139e-10, 1.406804e-10, 
    -1.13377e-10, 2.665999e-10, 2.864553e-10, -6.085799e-11, 9.011814e-11, 
    -5.342642e-10, 5.125909e-10, 2.027711e-11, 1.007416e-10, -4.890879e-10, 
    -8.128254e-10, -4.615472e-10, 1.60059e-09, 2.237122e-09, 1.326079e-09, 
    -1.027374e-10, -2.594973e-10, 5.14504e-11, -3.387086e-10, -2.060645e-10, 
    1.769251e-11, 1.758949e-11, -2.229328e-13, -8.508749e-12, -3.428369e-11,
  -2.325784e-10, 1.451578e-09, 2.516895e-09, 2.55579e-09, -7.532499e-10, 
    -3.626646e-10, 7.141772e-10, -5.312621e-10, 1.467594e-09, -2.032614e-10, 
    -1.031896e-09, 8.369447e-10, -1.952206e-09, -3.034764e-10, -3.994423e-10, 
    -2.922199e-10, -1.15353e-09, 8.506973e-11, -4.090772e-11, 9.762502e-11, 
    2.020037e-10, -7.805312e-12, 8.553158e-11, 1.58111e-09, -5.87524e-09, 
    4.682331e-09, 4.690399e-10, -3.643553e-09, -1.62192e-10, 1.447955e-09, 
    2.887287e-09, -9.842331e-10, -1.70451e-09, 8.541829e-09, 1.340901e-10, 
    1.101369e-08, -6.885514e-11, 9.510615e-12, -3.972421e-09, 1.763546e-10, 
    8.011369e-12, -1.809362e-10, 3.8618e-11, -4.880187e-10, -6.201795e-10, 
    3.411422e-10, 2.331468e-10, 1.020922e-09, -2.981302e-10, 1.870868e-10, 
    5.249525e-10, -8.446257e-10, -2.752001e-11, 3.381949e-10, 2.918519e-11, 
    5.27578e-12, 2.307583e-09, -4.498233e-11, -2.896118e-09, -2.135982e-09, 
    -2.713172e-10, -2.360174e-10, -1.261817e-10, 7.617799e-11, -3.245262e-11, 
    9.174254e-09, -1.48842e-09, 1.450854e-09, 1.908216e-09, -9.872636e-11, 
    1.119798e-09, 1.850534e-09, -2.768026e-10, -1.563979e-09, -2.128694e-10, 
    3.674572e-11, 8.011369e-13, 8.958878e-11, -1.185256e-11, 4.738148e-10, 
    1.014691e-10, 1.630809e-09, -7.448264e-11, 3.905807e-09, -3.458428e-09, 
    1.304695e-09, 3.002352e-09, 1.534417e-11, 1.732768e-09, 5.68722e-10, 
    -3.443294e-09, -2.488129e-10, 3.666401e-12, -1.471904e-09, 8.182859e-10, 
    -1.079421e-10, 5.256133e-10, 8.31843e-10, -2.254588e-10, 1.69748e-10, 
    -1.120075e-09, 4.298064e-10, 7.179146e-12, 1.086544e-10, -1.204061e-09, 
    -9.144294e-10, -5.685798e-10, 9.056684e-10, 1.968612e-09, 2.718632e-09, 
    -5.811174e-11, -5.431566e-10, -8.629186e-11, 2.725287e-11, -3.82304e-10, 
    3.025136e-11, 2.447642e-11, 2.01883e-12, -8.949286e-12, -8.185808e-11,
  4.640874e-10, 2.100723e-09, 4.795488e-10, -6.667413e-10, -3.579242e-09, 
    -6.955894e-10, -1.014978e-09, 5.861871e-10, 9.97364e-10, 6.395489e-10, 
    -7.900915e-10, 2.871477e-09, -3.393151e-09, -1.956941e-10, -1.484288e-10, 
    -5.815515e-10, -2.789493e-09, 5.107736e-11, -4.304823e-11, 1.170015e-10, 
    2.766605e-10, 5.157474e-11, 9.496404e-12, 1.214691e-09, -2.523954e-10, 
    5.016805e-09, 6.883347e-10, -5.91367e-10, -1.225725e-09, -4.220677e-09, 
    1.339022e-08, 1.091145e-10, 9.265939e-10, 7.379217e-09, 2.195755e-10, 
    1.680704e-08, -3.038871e-10, 1.210054e-11, -4.948799e-09, 2.510866e-10, 
    -3.263023e-11, -4.304148e-10, -2.34003e-10, -1.819349e-10, -6.355627e-10, 
    2.874145e-12, 8.131096e-11, 1.317211e-09, -2.560391e-10, 3.7618e-10, 
    4.370033e-10, -1.130569e-09, -3.323287e-10, 3.538282e-10, 7.389644e-12, 
    7.506884e-12, 2.861203e-09, -6.880256e-11, -2.529225e-09, -1.025507e-09, 
    -1.759979e-10, -2.356551e-10, -1.110401e-10, 5.979366e-10, -1.170768e-10, 
    2.073807e-08, -1.143615e-09, 4.294272e-10, 7.681809e-09, 7.170264e-10, 
    -5.940954e-10, 1.460084e-09, -3.238192e-10, -7.687468e-10, 6.797549e-11, 
    8.596501e-11, -3.165468e-12, 1.070184e-10, -1.414925e-10, 1.239364e-10, 
    3.445884e-10, 2.510834e-09, -5.682566e-11, 6.955336e-09, 1.695003e-09, 
    1.011138e-10, 3.692296e-09, 4.675726e-11, 1.697938e-09, 2.160938e-10, 
    -4.086825e-09, 4.282107e-10, -2.462031e-12, -1.138132e-08, 1.336961e-09, 
    -9.8661e-11, 5.048953e-10, 2.306397e-09, -4.136034e-10, 1.465402e-10, 
    -1.999734e-09, 4.982974e-10, -3.629097e-12, 8.447465e-11, -1.62208e-09, 
    -4.789165e-10, -8.355379e-10, 5.973426e-10, 3.005542e-09, 4.643955e-09, 
    2.234408e-10, -6.875602e-10, -1.622702e-10, -1.159545e-09, -6.494609e-10, 
    4.099903e-11, 3.282352e-11, 2.346701e-11, -2.701128e-11, -9.78666e-11,
  1.898144e-09, 6.299246e-09, 1.355858e-09, -1.580764e-08, -2.490935e-09, 
    3.733504e-09, -6.442974e-09, 2.148539e-09, -5.670984e-10, 1.148209e-09, 
    -4.849596e-10, 2.149164e-09, -2.214307e-09, 7.379413e-10, -6.493508e-10, 
    -1.126813e-09, -3.541075e-09, -4.558274e-10, 1.982414e-11, 1.510614e-10, 
    3.575735e-10, 1.465423e-10, 1.915623e-11, 1.32593e-09, 3.362743e-09, 
    1.606026e-09, -1.750152e-09, 2.359798e-09, -7.603916e-09, -6.192948e-09, 
    1.966919e-08, 2.014048e-09, 1.956266e-10, 4.293554e-09, 8.989787e-11, 
    2.62296e-08, -5.165248e-10, 1.591616e-11, -1.092454e-08, 1.833968e-10, 
    6.246239e-10, -7.525216e-10, -4.234479e-10, -2.169029e-10, -2.600615e-09, 
    -1.434074e-09, -2.553122e-10, 2.004391e-09, 2.984507e-10, 1.779359e-10, 
    4.852936e-10, -6.90477e-10, -2.955147e-10, 3.392529e-10, 5.193854e-11, 
    -1.11271e-11, 3.586337e-09, -1.112312e-10, -6.537277e-10, 1.913147e-09, 
    -1.609237e-10, -3.126956e-10, -3.00787e-10, 1.504606e-09, -1.181297e-09, 
    2.136886e-08, -8.175789e-10, -2.938748e-09, 4.169181e-09, -1.266187e-10, 
    -2.346923e-09, 2.545733e-10, -2.111449e-10, 2.934968e-09, 1.916109e-09, 
    1.742535e-10, -2.462741e-11, 1.548059e-10, -2.631111e-10, -1.172026e-09, 
    7.707541e-10, 3.52473e-09, 4.249046e-12, 8.672515e-09, 4.398004e-09, 
    2.2834e-10, 2.871957e-09, 7.935341e-11, 1.579796e-09, -1.287503e-11, 
    -5.47459e-09, 6.292e-11, -1.155342e-11, -2.326264e-08, 1.546709e-10, 
    -1.774936e-11, -1.113335e-10, 3.430813e-09, -5.040874e-10, 9.038104e-11, 
    -2.831797e-09, 7.962004e-10, -2.251355e-11, 4.933476e-11, 1.420801e-10, 
    6.157848e-10, -1.137096e-09, 4.488356e-10, 1.638796e-09, 6.173792e-09, 
    4.536957e-10, -6.542962e-10, -2.745537e-11, -1.08588e-09, -8.276402e-10, 
    5.96259e-11, 4.13003e-11, 6.687007e-11, -6.652279e-11, -1.386127e-10,
  2.979959e-09, 9.244474e-09, 9.119503e-09, -1.383057e-09, 2.038888e-09, 
    -4.21673e-09, -8.62164e-09, 7.328822e-10, 3.467733e-10, 4.193623e-10, 
    1.645702e-09, -9.916334e-10, -2.417494e-09, 1.544322e-09, -1.280199e-09, 
    -1.344205e-10, -4.464713e-09, -2.018652e-09, -1.999823e-11, 
    -1.019487e-10, 5.560707e-10, 2.730758e-10, 5.684342e-12, 7.523511e-10, 
    3.524264e-09, -1.601876e-09, -2.515208e-09, -1.172921e-08, -2.455124e-09, 
    -1.303601e-08, 2.669537e-09, -4.309982e-09, -4.097217e-09, 2.640434e-09, 
    -1.720082e-10, 3.711904e-08, -8.347513e-10, 3.241851e-11, -4.456069e-09, 
    -5.568211e-10, 8.369057e-10, -1.049699e-09, -1.704024e-10, -4.864416e-10, 
    -5.868685e-09, -2.005237e-09, -5.297096e-10, 2.379707e-09, 1.390674e-09, 
    1.276224e-10, 7.204832e-10, 5.921663e-10, -4.190355e-10, 4.309129e-10, 
    1.530864e-10, -6.579626e-11, 4.352302e-09, -1.692598e-10, 7.57052e-10, 
    1.448682e-08, -4.169465e-10, -5.279333e-10, -3.792024e-10, 1.580338e-09, 
    -2.705236e-10, 1.607248e-08, -2.666894e-09, -4.209738e-09, 4.580301e-09, 
    -1.984489e-09, -1.992589e-09, 4.317513e-09, -2.676728e-09, 9.485461e-10, 
    4.395556e-09, 2.125091e-10, -4.571987e-11, 2.49166e-10, -3.456648e-10, 
    -1.310895e-09, 1.500055e-09, 4.266689e-09, 9.755752e-11, 9.619328e-09, 
    2.806814e-09, 1.21679e-09, 9.670771e-10, 1.844569e-10, 1.63987e-09, 
    4.246203e-11, -1.794831e-10, -3.179308e-10, -2.653877e-11, -2.709577e-08, 
    -2.19103e-10, 1.101046e-09, -1.195878e-09, 2.298975e-09, -4.683613e-10, 
    5.682068e-11, -2.189779e-09, 1.548777e-09, -8.279244e-11, 2.170708e-12, 
    5.697132e-10, 6.924665e-10, 9.657981e-10, 2.490907e-09, 1.910337e-09, 
    6.507207e-09, 4.705782e-10, -6.130563e-10, 1.054445e-10, -1.721503e-10, 
    -1.023807e-09, 9.091253e-11, 5.617196e-11, 1.163007e-10, -9.717027e-11, 
    -2.612524e-10,
  2.858968e-09, 8.63858e-09, 5.456428e-09, 1.770655e-08, 3.017902e-09, 
    -6.20048e-10, -2.470614e-09, -4.62785e-09, 4.201155e-09, -3.426806e-10, 
    2.135721e-09, -3.021512e-09, -2.389868e-09, 4.226706e-09, 5.592824e-10, 
    8.828978e-10, -7.263623e-09, -2.012584e-09, -2.986447e-10, -4.835954e-10, 
    7.202914e-10, 6.916707e-10, -1.536193e-10, 3.897469e-10, 2.489429e-09, 
    2.315232e-10, -1.779767e-10, -1.541122e-08, 1.132807e-08, -2.003449e-08, 
    -7.456691e-09, -5.569376e-09, -9.477873e-09, 2.956199e-09, -1.644764e-10, 
    4.391364e-08, -1.244925e-09, 6.595258e-11, -1.526871e-08, -1.681721e-09, 
    6.349641e-10, -1.564814e-09, 4.366996e-11, -8.584529e-10, -1.276666e-08, 
    3.060222e-09, -5.59524e-10, 2.751975e-09, 2.498143e-09, 9.69127e-11, 
    1.132857e-09, 1.369642e-09, -7.427615e-10, 6.373e-10, 1.832312e-10, 
    -1.34122e-10, 5.297096e-09, -3.135852e-10, -6.74703e-10, 1.639494e-08, 
    -9.14838e-10, -5.427978e-10, -1.47196e-10, 5.839922e-10, 1.07496e-09, 
    1.329184e-08, -4.598121e-09, -2.056055e-09, 4.154458e-09, -5.120938e-09, 
    -6.139658e-10, 3.791192e-08, -4.448765e-09, -4.103015e-09, 6.651646e-09, 
    1.239755e-10, -6.420819e-11, 4.910987e-10, -4.097451e-10, 4.030483e-10, 
    3.007784e-09, 5.733807e-09, 1.737703e-10, 9.319479e-09, -1.484807e-09, 
    2.613888e-09, -2.750539e-09, 3.8591e-10, 1.774598e-09, 9.894165e-10, 
    1.080136e-08, -1.228107e-09, 2.846434e-11, -1.807908e-08, -3.038281e-10, 
    2.917153e-09, -1.85845e-09, -6.41478e-10, -4.97721e-10, -2.962679e-11, 
    -1.810378e-09, 2.317483e-09, -1.644924e-10, -8.683543e-11, 5.712764e-10, 
    9.729035e-10, 2.896087e-09, 2.317989e-09, 1.285883e-09, 8.073641e-09, 
    1.594174e-09, -5.064749e-10, -2.842455e-10, -1.546198e-09, -1.448541e-09, 
    4.289973e-11, 9.790924e-11, 9.523049e-11, -9.951862e-11, -4.115748e-10,
  2.412719e-09, 6.027335e-09, -4.18936e-10, 3.938396e-09, 8.964776e-10, 
    -1.571721e-10, -3.275886e-10, -1.333461e-08, 3.561922e-09, -2.5085e-10, 
    1.382318e-09, -1.330932e-09, -1.431658e-09, 1.267551e-09, 4.03935e-09, 
    1.854295e-09, -5.106415e-09, -7.437961e-10, -4.718927e-10, -1.147669e-10, 
    1.293301e-09, 7.556764e-10, -1.074341e-10, 1.607532e-10, 5.233005e-10, 
    2.978538e-09, -3.295327e-09, -1.384268e-08, 1.284809e-08, -1.786611e-08, 
    2.034142e-09, -7.035851e-09, -1.143786e-08, 2.920444e-09, 1.078888e-10, 
    5.060082e-08, -1.273679e-09, 7.349854e-11, -4.153219e-08, -2.989015e-09, 
    1.275122e-10, -2.36264e-09, -2.164882e-10, -1.483866e-09, -1.554042e-08, 
    9.12928e-09, -2.499519e-09, 2.434589e-09, 2.996546e-09, 7.16085e-11, 
    1.658897e-09, 4.260983e-10, -5.89199e-10, 9.534119e-10, 1.011628e-10, 
    -1.066667e-10, 5.481184e-09, 9.806056e-11, -5.124031e-09, 8.108863e-09, 
    -1.656872e-09, -1.897433e-10, -4.718004e-12, 1.217779e-09, 1.283036e-09, 
    3.587047e-09, -5.780407e-09, -4.06709e-09, 6.012272e-09, -4.203685e-09, 
    3.634e-10, 3.760283e-08, -3.122125e-09, 2.591946e-09, 6.59349e-09, 
    -2.216893e-12, -6.426149e-11, 6.311041e-10, -4.841368e-10, -4.197886e-10, 
    4.835073e-09, 8.034594e-09, 2.317222e-10, 6.86839e-09, -5.502784e-09, 
    2.885315e-09, -7.80534e-09, 5.154561e-10, 2.41381e-09, 2.473314e-09, 
    1.177727e-08, -2.480419e-09, 2.455351e-10, -1.0684e-08, -2.891852e-09, 
    6.12812e-10, -2.607919e-09, -4.975391e-09, -1.105263e-09, -1.797048e-10, 
    -1.13306e-09, 2.253099e-09, -1.601386e-10, -1.268923e-10, 9.82368e-10, 
    8.652705e-10, 1.688761e-09, 2.449212e-09, 4.227445e-10, 1.000234e-08, 
    3.803393e-09, -1.503508e-10, -2.102865e-09, -4.958224e-09, -2.25009e-09, 
    -5.534844e-11, 1.848406e-10, -1.731948e-11, -8.851941e-11, -4.662297e-10,
  2.083652e-09, 3.883031e-09, -1.47071e-09, 2.567674e-09, 4.65036e-10, 
    -6.471623e-10, 7.09349e-10, -1.429368e-08, 1.082128e-09, 3.279808e-09, 
    9.079031e-10, -1.451554e-09, -1.505555e-09, -6.681603e-09, 2.004867e-09, 
    -1.616769e-09, 1.684344e-09, 1.102393e-09, -9.687398e-10, 8.020038e-10, 
    3.067839e-09, 1.10748e-09, 5.545644e-10, 5.23471e-10, -1.158242e-09, 
    1.212356e-09, -2.559261e-09, -2.296866e-08, 2.426702e-09, -3.960281e-10, 
    2.539252e-09, -9.359439e-09, -1.522397e-08, 2.195691e-09, 8.782308e-11, 
    5.854486e-08, -1.786782e-09, 5.586287e-11, -5.672405e-08, -5.087776e-09, 
    4.946844e-09, -2.188131e-09, -6.290577e-10, -1.996765e-09, -6.03535e-09, 
    1.396637e-08, -9.380329e-09, 1.608825e-09, 2.728041e-09, 8.076029e-11, 
    1.925905e-09, -1.433591e-10, -1.002376e-10, 1.307774e-09, 5.054076e-10, 
    2.02931e-11, 3.078071e-09, 1.655201e-09, -1.159638e-08, 2.708695e-09, 
    -4.637741e-09, 1.756462e-10, -8.930101e-10, 2.19751e-09, -8.377015e-10, 
    1.731848e-08, -6.346454e-09, -1.289811e-08, 3.753996e-09, -6.436323e-09, 
    -8.907364e-11, 3.142412e-08, -9.455903e-10, 7.724282e-09, 3.873486e-09, 
    -1.284661e-10, -1.673328e-11, 5.941985e-10, -6.292396e-10, 2.470074e-09, 
    6.802054e-09, 1.020948e-08, 2.14925e-10, 2.912657e-10, -2.407035e-09, 
    1.51482e-09, -4.674803e-09, 6.397727e-10, 4.342705e-09, 4.838e-09, 
    9.470341e-09, -7.659684e-09, 6.701839e-10, -1.258875e-08, -1.959052e-09, 
    -1.513271e-08, 6.408754e-10, -4.829928e-09, -2.054662e-09, -3.433001e-10, 
    3.738592e-10, 1.044032e-09, -1.636487e-10, -1.933032e-11, 2.286072e-09, 
    -2.735874e-10, 1.366914e-09, 1.709736e-09, -4.141327e-09, 1.179831e-08, 
    3.977163e-09, -1.742819e-10, -4.63308e-09, -8.605696e-09, -1.849344e-09, 
    -6.663185e-11, 3.395826e-10, -4.193801e-11, -7.509371e-11, -7.41295e-10,
  6.533583e-10, -6.772325e-10, -1.448086e-09, 1.458091e-09, 1.023238e-09, 
    5.478569e-10, 9.003998e-11, -4.782294e-09, -3.740013e-09, 5.741072e-09, 
    2.052843e-09, -2.806189e-09, -3.391563e-09, -5.696506e-09, -1.208565e-08, 
    -3.97614e-09, 6.055314e-09, 3.353705e-09, -2.770236e-09, 1.46548e-09, 
    3.998593e-09, 2.093941e-09, 1.348724e-09, 9.015366e-10, -2.303864e-10, 
    -8.683969e-10, 6.356686e-09, -1.492384e-08, -2.484057e-11, -3.822265e-09, 
    2.696538e-09, -1.078757e-08, -2.242621e-08, 2.259924e-09, -1.660453e-09, 
    6.040966e-08, -1.717558e-09, 8.036238e-11, -3.740257e-08, -9.575712e-09, 
    1.540503e-09, 6.090772e-10, -7.99389e-10, -1.941065e-09, -9.746827e-09, 
    1.709168e-08, -2.236007e-08, -1.57641e-10, 2.226886e-09, 3.252154e-11, 
    1.213316e-09, 1.074511e-09, 1.943982e-09, 1.791807e-09, 1.343713e-09, 
    1.186606e-10, -2.800448e-09, 3.634051e-09, -1.596353e-08, -6.536801e-09, 
    -1.172685e-08, -6.474465e-11, -1.862986e-09, 2.400384e-09, -6.330776e-09, 
    3.0553e-08, -4.283436e-09, -2.847679e-08, 1.09539e-08, -7.395158e-09, 
    -9.926566e-10, 6.193716e-09, -2.157776e-10, 5.816617e-09, 1.931011e-09, 
    -1.668923e-10, -2.280842e-12, 4.473861e-10, -8.648243e-10, 8.031179e-09, 
    9.980198e-09, 1.036265e-08, 3.546177e-10, -2.477293e-09, 2.842398e-09, 
    1.150568e-09, 1.434444e-09, 9.251835e-10, 9.168332e-09, 9.296997e-09, 
    9.970506e-09, -1.454646e-08, 1.096211e-09, -1.875628e-08, -1.103729e-09, 
    -2.307624e-08, 1.98371e-09, 6.431719e-09, -2.805848e-09, -4.373192e-10, 
    -4.845901e-10, 6.456702e-11, -6.889529e-10, 3.002292e-10, 3.774062e-09, 
    -6.944504e-09, 1.985313e-09, -2.091724e-09, -1.259764e-09, 1.1569e-08, 
    1.770957e-09, -2.392539e-10, -8.646623e-09, -1.317812e-08, -1.046033e-09, 
    -6.118626e-11, 4.962928e-10, -1.249063e-10, -4.723333e-11, -4.354206e-10,
  -9.013092e-10, -5.043034e-09, -2.99832e-09, -3.858531e-10, 8.4151e-10, 
    2.21678e-09, -7.77618e-11, 4.440949e-09, -1.100472e-08, 2.513559e-09, 
    5.772904e-09, -6.688197e-10, -2.774073e-09, 1.812339e-09, -1.436422e-08, 
    -4.958042e-09, 1.050517e-08, 5.49619e-09, -5.747196e-09, 1.364754e-09, 
    2.815341e-09, 2.398224e-10, 2.083141e-09, 2.027946e-09, 2.200409e-10, 
    -1.464571e-09, -1.322712e-08, -2.315278e-08, -1.25911e-08, -9.143946e-09, 
    -2.320292e-09, -1.098164e-08, -2.988133e-08, 1.804665e-09, -4.571291e-09, 
    5.914984e-08, -1.286583e-09, 1.118394e-10, -2.227847e-08, -1.589465e-08, 
    5.357833e-09, 4.061974e-09, -5.364171e-10, -1.89499e-09, -2.016247e-08, 
    1.962388e-08, -2.989614e-08, -4.196721e-09, 1.114915e-09, 1.715605e-11, 
    -7.081695e-10, 2.614399e-09, 3.882451e-09, 2.37909e-09, 2.318154e-09, 
    1.812168e-10, -8.612403e-09, 6.160104e-09, -2.124972e-08, -1.867571e-08, 
    -5.303889e-09, 2.210641e-10, -2.80528e-09, -3.661057e-10, -7.893209e-09, 
    2.665712e-08, 1.494698e-09, -3.999958e-08, 1.436399e-08, -2.347747e-09, 
    -1.030514e-09, -1.936155e-08, -8.804818e-09, 6.822347e-10, 2.534586e-09, 
    -1.677449e-10, -7.934631e-11, 5.62153e-10, -1.132197e-09, 1.074596e-08, 
    1.513078e-08, 9.896517e-09, 6.134258e-10, -3.673335e-09, 5.975039e-09, 
    1.576495e-09, 3.646846e-09, 8.581651e-10, 2.06536e-08, 1.638585e-08, 
    1.27302e-08, -1.918812e-08, 1.406463e-09, -3.63682e-08, 2.420961e-10, 
    -2.654506e-08, 2.686409e-09, 2.19145e-08, -4.790536e-09, -4.302933e-10, 
    -1.754984e-09, -5.064997e-10, -1.445105e-09, 9.787051e-10, 1.008817e-08, 
    3.168054e-09, 1.973888e-09, -4.770243e-09, 5.112554e-09, 7.450865e-09, 
    8.6402e-10, -2.052332e-09, -6.401763e-09, -2.555788e-08, -6.283699e-09, 
    -1.872991e-11, 6.394458e-10, -1.332605e-10, -4.942891e-11, -1.365379e-10,
  -1.613728e-09, -1.939441e-09, -2.139586e-09, -1.755325e-09, 2.549427e-10, 
    1.497312e-09, 8.654979e-10, 5.368292e-09, -1.589007e-08, -3.667481e-09, 
    3.099672e-09, -3.616776e-09, 4.368417e-10, 4.200331e-09, 3.183231e-09, 
    -5.785927e-09, 1.398085e-08, 6.855885e-09, -9.933117e-09, 1.454623e-10, 
    1.785224e-09, -2.843308e-10, 2.398224e-09, 3.170726e-09, 3.374225e-10, 
    -2.451657e-10, 3.326682e-08, -2.352027e-08, -5.48834e-08, -6.685184e-09, 
    1.160601e-08, -1.042503e-08, -3.200296e-08, 2.708703e-09, -3.005198e-09, 
    5.85128e-08, 7.553183e-10, 1.537686e-10, -1.184679e-08, -2.219388e-08, 
    1.590148e-08, 3.957268e-09, 4.011866e-10, -2.739885e-09, -1.491071e-08, 
    1.17862e-08, -2.150506e-08, -1.245726e-08, -6.994014e-10, 6.743051e-12, 
    -4.658126e-09, 5.310994e-09, 3.987753e-09, 3.153798e-09, 3.381422e-09, 
    1.77522e-10, -1.026234e-08, 1.432536e-08, -4.72804e-08, -1.17307e-08, 
    6.251412e-09, 1.474916e-09, -2.752245e-09, -6.169444e-09, 1.782041e-09, 
    9.802648e-09, 7.685571e-09, -3.870775e-08, 2.257264e-08, 7.628955e-10, 
    -1.562296e-08, -4.272692e-08, -2.086205e-08, -2.143963e-09, 5.594512e-09, 
    1.284661e-10, 2.647482e-11, 2.292353e-10, -1.437451e-09, 7.149424e-09, 
    2.307016e-08, 1.040504e-08, 1.020908e-09, -8.581651e-10, 1.169894e-09, 
    6.386358e-10, 3.285606e-09, 3.220748e-10, 4.391363e-08, 3.032824e-08, 
    9.855796e-09, -3.134984e-08, 1.393772e-09, -7.298311e-08, 4.331469e-11, 
    -1.829862e-08, -2.31346e-09, 2.949309e-08, -1.044208e-08, -3.802825e-10, 
    -2.988088e-09, -4.426397e-10, -2.053667e-09, 2.084178e-09, 6.131415e-09, 
    3.732737e-09, -1.793524e-09, -9.835048e-10, 5.068557e-09, 2.843763e-09, 
    -7.89953e-10, -3.15282e-09, 4.928097e-09, -3.482785e-08, -1.620742e-08, 
    4.095e-11, -9.029577e-11, -1.400089e-10, -4.640555e-11, 9.799237e-10,
  -2.770093e-09, -3.633431e-10, -2.282832e-10, -1.906699e-09, -2.361787e-09, 
    -1.831324e-09, -2.857917e-09, -1.571266e-09, -1.070202e-08, 
    -1.148794e-08, -3.942489e-09, -4.650815e-09, 6.667051e-09, 2.601496e-09, 
    1.037967e-08, -7.064091e-09, 1.796878e-08, 6.494162e-09, -1.414442e-08, 
    -8.94147e-10, 3.783441e-09, 3.541629e-09, -7.716494e-10, 3.969262e-09, 
    6.946266e-11, 7.246399e-10, 6.582951e-08, -1.668087e-08, -9.522444e-08, 
    -8.264465e-09, 1.032402e-08, -1.034419e-08, -3.058818e-08, 8.155041e-09, 
    3.82181e-09, 7.386808e-08, 3.252637e-09, 2.525624e-10, 1.920796e-09, 
    -3.335916e-08, 2.282755e-08, 4.010587e-09, 1.726235e-09, -6.69868e-09, 
    -3.294815e-09, -6.394373e-09, -2.50526e-09, -2.578879e-08, -8.007669e-09, 
    2.041389e-11, 3.44798e-10, 3.709999e-09, -2.021893e-08, 4.346839e-09, 
    4.423258e-09, 8.932943e-11, -6.782386e-09, 1.458756e-08, -6.023805e-08, 
    1.499546e-08, 8.265374e-09, 2.238721e-09, -3.390312e-09, -1.357435e-08, 
    7.923677e-09, 7.522601e-09, 7.872188e-09, -3.771112e-08, 4.116987e-08, 
    2.884235e-10, -5.279713e-08, -5.411061e-08, -2.090184e-08, -3.069431e-09, 
    9.337396e-09, 7.927952e-10, -1.370779e-10, -3.935554e-10, -1.995757e-09, 
    2.51714e-09, 3.243289e-08, 1.435269e-08, 1.542361e-09, 5.275069e-10, 
    1.121236e-09, -1.697231e-09, 5.356867e-09, 2.270951e-09, 7.106315e-08, 
    5.362475e-08, 2.878437e-09, -4.903559e-08, 8.843131e-10, -1.038481e-07, 
    -6.818937e-10, -3.892018e-09, -6.563187e-09, 1.774839e-08, -1.126239e-08, 
    -5.840093e-10, -2.728996e-09, 7.071961e-10, -3.267598e-09, 3.377284e-09, 
    1.348724e-09, -5.376762e-09, -4.39627e-09, 2.647425e-09, 1.893568e-09, 
    1.506919e-09, 2.302158e-11, -2.094055e-09, 1.485603e-09, -2.988469e-08, 
    -1.572198e-08, 1.395278e-10, -6.047784e-10, -1.615383e-10, -1.548628e-11, 
    2.217405e-09,
  -4.272295e-09, 9.549694e-12, -9.731593e-11, -1.139824e-09, -2.505772e-09, 
    -2.774186e-09, -9.152586e-09, -9.44533e-09, 4.830099e-09, -8.460063e-09, 
    -5.099366e-09, 1.472472e-09, 4.665139e-09, 3.670152e-09, 2.45447e-08, 
    -7.947586e-09, 1.948803e-08, 4.274341e-09, -1.623923e-08, 4.819753e-10, 
    5.97214e-09, 9.860685e-09, 7.416361e-10, 5.173206e-09, -5.79746e-10, 
    6.315304e-10, -1.991583e-08, -1.108464e-08, -6.079455e-08, -1.371149e-08, 
    8.951133e-10, -1.665018e-08, -3.369996e-08, 2.000269e-08, 8.647703e-09, 
    8.419607e-08, 5.785665e-09, 4.083702e-10, 1.16035e-08, -4.265874e-08, 
    3.387661e-08, 2.825175e-09, 4.306742e-09, -7.82723e-09, 3.483427e-08, 
    -7.234917e-09, 2.076814e-08, -4.492908e-08, -2.119473e-08, 9.778844e-11, 
    6.586873e-09, 1.174612e-09, -5.411098e-08, 6.292953e-09, 5.11611e-09, 
    2.268052e-11, 7.151186e-09, 2.450085e-08, -3.214633e-08, 3.356109e-08, 
    2.433353e-09, -1.808985e-09, -4.512174e-09, -1.711732e-08, 9.197243e-09, 
    -5.202139e-09, 2.306575e-08, -1.871848e-08, 6.648941e-08, 1.449962e-09, 
    -8.513581e-08, -2.071289e-08, -2.766251e-08, -4.305605e-09, 1.241784e-08, 
    1.482761e-09, -1.869509e-10, -1.912085e-09, -2.564388e-09, 3.400373e-10, 
    3.201799e-08, 2.681975e-08, 2.289426e-09, 1.111061e-09, -5.317702e-10, 
    -2.724221e-09, 4.170431e-09, 7.318988e-09, 8.692848e-08, 8.972896e-08, 
    2.142997e-11, -6.086109e-08, -8.341914e-10, -1.502193e-07, 1.327408e-09, 
    -2.359739e-08, -1.330246e-08, 1.396364e-08, -1.427566e-08, -1.486399e-09, 
    3.638547e-10, 4.735092e-10, -7.253004e-09, 5.02008e-09, 1.04535e-10, 
    -9.94703e-09, 3.495302e-09, 4.878245e-09, 5.190941e-10, 1.186834e-09, 
    8.306529e-10, -5.055085e-10, -3.069658e-09, -1.729359e-08, -9.720793e-10, 
    3.468642e-10, -8.808811e-10, -2.300915e-10, 3.932854e-11, 2.319041e-09,
  -2.879233e-09, -2.512479e-11, 2.383103e-09, 1.590934e-09, -1.352646e-09, 
    -1.596277e-09, -1.101967e-08, -1.230671e-08, 2.071533e-08, 2.049092e-09, 
    5.28496e-09, 7.357016e-09, 3.523155e-10, 1.386752e-09, 1.716217e-08, 
    -2.888942e-09, 2.098147e-08, 5.065885e-10, -1.767069e-08, 5.393531e-09, 
    1.675176e-09, 2.112643e-09, 2.916295e-09, 5.404559e-09, -8.300276e-10, 
    -1.27784e-09, 1.080025e-11, -2.926117e-08, -2.963475e-08, -1.148419e-08, 
    -2.710442e-08, -2.944705e-08, -4.682897e-08, 3.463867e-08, 9.797873e-09, 
    8.674408e-08, 6.999335e-09, 6.717187e-10, 1.8739e-09, -5.286191e-08, 
    5.664992e-08, 1.156081e-09, 8.610641e-09, 1.494286e-08, 2.328932e-08, 
    9.299333e-08, 3.914749e-08, -6.631043e-08, -3.82975e-08, 1.695071e-10, 
    1.391409e-08, 3.308855e-09, -5.150893e-08, 5.523998e-09, 5.874881e-09, 
    -1.758735e-10, 3.563844e-08, 2.669884e-08, -1.660086e-08, 2.381901e-08, 
    -4.004733e-09, -5.555421e-09, -2.979732e-09, -1.535e-08, 6.446634e-09, 
    -1.818808e-08, 1.430942e-08, -1.905562e-08, 3.88909e-08, 6.108621e-09, 
    -1.163905e-07, 7.329368e-08, -3.497485e-08, -8.298002e-10, 1.225172e-08, 
    2.29636e-09, -2.402061e-10, -3.809902e-09, -2.648378e-09, 3.308287e-10, 
    3.740558e-08, 4.309647e-08, 3.293962e-09, -2.975185e-10, -4.738013e-09, 
    3.943228e-09, -8.537882e-10, 8.3553e-09, 8.358792e-08, 1.300481e-07, 
    -3.551804e-09, -6.260391e-08, -2.590781e-09, -1.881854e-07, 
    -1.468266e-08, -7.203054e-08, -2.363693e-08, 3.700882e-08, -1.35384e-08, 
    -3.422951e-09, 3.00065e-09, 1.19698e-10, -1.517434e-08, 5.037812e-09, 
    -2.768502e-09, -1.100034e-08, -2.166416e-09, 4.374328e-09, 4.081357e-10, 
    7.12248e-10, 4.891945e-10, -4.102958e-10, -3.292826e-09, -4.207095e-09, 
    1.358785e-08, 4.016329e-10, -7.625118e-10, -1.416502e-10, 1.031353e-10, 
    3.050673e-09,
  -2.172612e-09, -5.690026e-11, 2.243326e-09, 2.027747e-08, 1.211276e-09, 
    -8.429311e-10, -8.82693e-09, -7.918004e-09, 1.823395e-08, 1.847064e-08, 
    1.636869e-08, 3.970229e-09, -1.073374e-09, -7.414087e-10, -1.0603e-09, 
    1.403965e-08, 1.840843e-08, 3.4089e-10, -2.075724e-08, 1.216875e-08, 
    -1.694212e-08, -4.491034e-08, -3.302324e-08, -2.726495e-09, 1.156025e-09, 
    -4.992955e-09, -2.117417e-10, -3.660858e-08, -2.239523e-08, 2.342705e-08, 
    -6.829549e-08, -3.952204e-08, -7.062289e-08, 1.421898e-08, 1.59817e-08, 
    9.257752e-08, 7.249969e-09, 8.842846e-10, 6.954508e-09, -6.507346e-08, 
    8.162641e-08, 2.357012e-09, 1.222998e-08, 1.97644e-08, 1.40389e-08, 
    3.030726e-08, 4.606659e-08, -8.857802e-08, -5.568301e-08, 1.551044e-10, 
    8.580315e-09, -1.818233e-08, -6.503205e-09, 5.252389e-09, 6.646712e-09, 
    -3.22359e-10, 7.394334e-08, 3.998348e-08, -3.071776e-08, 1.087822e-08, 
    1.287901e-09, -4.253764e-09, 1.052172e-10, -1.399213e-08, 2.15058e-09, 
    -1.150676e-08, -5.50591e-09, 1.645009e-07, 2.771174e-09, 6.93143e-09, 
    -1.340118e-07, 5.708358e-08, -1.978827e-08, 3.532762e-09, 7.973267e-09, 
    3.359617e-09, -4.268941e-10, -6.583804e-09, -2.548816e-09, -2.268052e-11, 
    5.014317e-08, 4.345473e-08, 4.230742e-09, -3.518437e-09, -5.326228e-11, 
    7.995197e-09, 8.553172e-09, 5.948493e-09, 6.557748e-08, 1.468012e-07, 
    -6.77818e-09, -5.759602e-08, -3.093248e-09, -2.055027e-07, -2.640326e-08, 
    -1.284834e-07, -3.66099e-08, 5.031796e-08, -1.26484e-08, -6.045081e-09, 
    -1.631975e-10, -1.295213e-09, -2.589719e-08, 3.54661e-09, -2.29835e-09, 
    -1.729876e-08, -1.177756e-08, 1.357438e-08, 3.499906e-09, 1.330648e-09, 
    1.001865e-09, 6.17888e-11, -1.375099e-09, 5.853678e-09, 1.06981e-08, 
    6.410005e-10, -6.663896e-10, -1.352483e-10, 1.529017e-10, 5.248864e-09,
  5.763923e-10, -1.919034e-10, 1.207468e-09, 4.562673e-08, 5.077936e-09, 
    8.971483e-09, -7.820404e-09, -2.712454e-09, 3.340915e-09, 2.125887e-08, 
    1.552564e-08, -4.562253e-10, -1.904482e-09, -4.816343e-09, -2.380375e-09, 
    3.806554e-08, 4.772268e-09, 3.030152e-09, -2.511307e-08, 1.614023e-08, 
    -4.803951e-08, -3.96459e-08, -3.881166e-08, -1.41182e-08, 3.003379e-09, 
    -5.714583e-09, 2.403056e-08, -3.108437e-08, -9.251949e-09, 4.230037e-08, 
    -7.98774e-08, 5.238576e-09, -8.673976e-08, -1.139597e-08, 1.888884e-08, 
    7.787196e-08, 8.340669e-09, 7.912746e-10, -1.601506e-09, -8.214386e-08, 
    1.041785e-07, 3.099785e-09, 1.051052e-08, 1.741542e-08, 1.612909e-08, 
    -1.431169e-08, 4.136592e-08, -1.142772e-07, -7.434687e-08, -1.462297e-10, 
    7.568289e-09, -4.511492e-08, 3.781017e-08, 9.245809e-09, 6.509418e-09, 
    -2.754632e-10, 1.006816e-07, 4.508986e-08, 2.942784e-10, 1.092019e-09, 
    9.225573e-09, -9.324594e-10, 1.000558e-09, -1.983738e-08, -6.663457e-09, 
    -4.465619e-08, -1.080241e-08, 1.616647e-07, -9.430778e-09, -2.435411e-08, 
    -1.29514e-07, -4.602839e-09, -3.978357e-09, 2.138108e-09, -9.18377e-09, 
    3.259061e-09, -7.356533e-10, -7.919681e-09, -2.079418e-09, 6.240271e-10, 
    5.607365e-08, 1.772155e-08, 4.307935e-09, -5.828042e-09, 5.01359e-09, 
    9.370751e-09, 3.218577e-08, 2.77123e-09, 4.424549e-08, 1.337704e-07, 
    -7.42682e-09, -4.76957e-08, -2.379835e-09, -1.506447e-07, -2.766137e-08, 
    -9.754096e-08, -5.416025e-08, 2.364357e-07, -8.8462e-09, -8.561165e-09, 
    -9.246833e-09, -6.443265e-09, -3.039307e-08, 3.159855e-09, -3.304763e-09, 
    -4.007029e-08, -1.911587e-08, 1.98329e-08, 1.007356e-08, 2.430397e-09, 
    1.885041e-09, 8.003553e-10, -1.236913e-10, 8.872803e-09, 9.723635e-10, 
    1.041519e-09, -6.680239e-10, -1.475904e-10, 2.234586e-10, 9.250471e-09,
  3.496211e-08, -1.076614e-10, 1.014882e-09, 4.512299e-08, 8.75923e-09, 
    2.970648e-08, -3.197101e-09, -4.569642e-09, -2.473598e-09, 4.357616e-10, 
    5.482093e-09, -3.222794e-09, -6.274377e-10, -3.11602e-08, -3.701643e-10, 
    4.432813e-08, -5.386461e-09, 2.310912e-09, -2.791943e-08, 1.274395e-08, 
    -6.493804e-08, -1.803642e-08, -1.09286e-08, -9.982045e-09, 4.82828e-09, 
    1.031708e-09, 5.518709e-07, -2.790944e-08, 1.244803e-08, 8.041184e-09, 
    -2.96767e-08, 1.765469e-07, -4.578158e-08, -2.759009e-08, 5.101811e-09, 
    4.818605e-08, 7.226459e-09, 6.045582e-10, 7.471385e-09, -1.036817e-07, 
    1.103418e-07, 1.515104e-09, 6.319453e-09, 1.544225e-08, 2.631737e-08, 
    -2.667264e-08, 2.956642e-08, -1.31541e-07, -7.6011e-08, -5.069225e-10, 
    -4.260713e-09, -5.343441e-08, 7.245798e-08, 1.543306e-08, 5.352905e-09, 
    -1.470539e-10, 9.852363e-08, 5.293507e-08, 6.249574e-08, -2.653749e-09, 
    6.327355e-09, -1.163016e-10, 1.606509e-09, -2.95146e-08, -1.86307e-08, 
    -5.452728e-08, -2.170339e-08, 7.791186e-08, 3.413447e-08, -4.616118e-08, 
    -1.040986e-07, -6.100379e-08, -1.122953e-08, 1.261128e-09, -3.486837e-08, 
    -1.548756e-09, -8.768524e-10, -8.610016e-09, -8.888037e-10, 2.231673e-10, 
    6.013488e-08, -2.762019e-09, 3.245816e-09, -5.946163e-09, 2.111619e-09, 
    -1.123919e-08, 1.915521e-08, -7.069048e-10, 2.616008e-08, 1.030975e-07, 
    -3.967671e-09, -3.160164e-08, -1.280341e-09, -3.504549e-08, 
    -2.903869e-08, -8.71234e-08, -8.105238e-08, 1.682123e-07, -3.432547e-09, 
    -1.060894e-08, -5.013158e-08, -1.246976e-08, -2.913952e-08, 2.380297e-09, 
    -1.508602e-08, -6.330583e-08, -3.411833e-08, 3.276011e-08, 1.83129e-08, 
    1.786475e-09, 3.227569e-10, 3.985861e-10, -1.21247e-09, 2.814886e-09, 
    -1.503281e-09, 1.47819e-09, -5.121876e-10, -2.459011e-10, 2.67562e-10, 
    1.84732e-08,
  3.66407e-08, 8.867573e-12, -9.987389e-10, 7.053359e-09, 5.618745e-09, 
    4.307935e-08, 6.881123e-09, -4.243816e-09, 1.41938e-09, -2.216666e-09, 
    -6.715595e-09, -1.076876e-08, 4.738467e-10, -5.842742e-08, -2.94574e-09, 
    2.979413e-08, -1.66009e-08, 2.489685e-09, -1.900793e-08, 5.983679e-09, 
    -4.262199e-08, -1.277783e-08, 8.118946e-09, -2.594561e-09, -3.981881e-09, 
    3.996433e-09, -1.585889e-07, -1.469971e-08, 7.467975e-09, -6.348091e-08, 
    -7.687049e-09, 2.298568e-07, 7.700351e-09, -6.058247e-08, -2.209606e-08, 
    3.516902e-08, 7.511494e-09, 3.622915e-10, 1.613103e-08, -1.228702e-07, 
    9.367191e-08, 1.263061e-09, -1.195161e-09, 9.476057e-09, 2.806325e-08, 
    -3.190917e-08, 1.641263e-08, -1.327105e-07, -5.960417e-08, -3.447823e-09, 
    -1.977757e-08, -6.674497e-08, 8.673078e-08, 1.969581e-08, 1.454347e-09, 
    -6.45116e-10, 9.255348e-08, 6.428951e-08, 1.075238e-07, -5.401745e-09, 
    2.230991e-09, -3.248033e-10, 2.442448e-09, -2.611068e-08, -3.147379e-08, 
    -3.964385e-08, -4.428523e-08, -3.624825e-08, 8.021163e-08, -2.089382e-08, 
    -1.086906e-07, -1.110116e-07, -9.503538e-09, 4.91741e-09, -4.433791e-08, 
    -1.444573e-08, 2.889919e-10, -1.139986e-08, 6.361347e-10, -5.325808e-08, 
    6.235865e-08, 2.239794e-08, 2.218314e-09, -4.701292e-09, -7.477752e-09, 
    -3.000491e-08, -5.4456e-11, -1.028866e-10, 1.606921e-08, 6.927712e-08, 
    1.05922e-09, -1.530575e-08, -1.375611e-11, 4.489655e-08, -1.182229e-08, 
    -2.021574e-08, -1.193435e-07, 4.566232e-09, -2.649585e-09, -1.304522e-08, 
    -5.991944e-08, -2.515635e-08, -2.013751e-08, 1.750038e-09, -6.890377e-08, 
    -5.417053e-08, -2.70129e-08, 3.387152e-08, 2.721674e-08, -1.666649e-10, 
    -3.734158e-09, -3.529976e-10, -2.803176e-09, -6.248001e-09, 3.933565e-11, 
    1.413264e-09, -8.861889e-11, -2.737224e-10, 2.677112e-10, 3.10738e-08,
  2.146959e-08, -1.689955e-10, -9.288158e-09, -3.190956e-08, 4.893025e-09, 
    3.944893e-08, 8.024188e-09, -5.492609e-09, -5.192476e-09, -3.907928e-09, 
    -2.265381e-09, -1.029895e-08, 4.874323e-10, -4.464783e-08, -1.181974e-08, 
    3.581768e-08, -2.470005e-08, 1.159265e-09, -1.839595e-10, -1.343039e-09, 
    1.291198e-09, -3.083568e-08, 7.450751e-09, -5.571962e-09, -1.136499e-08, 
    6.965024e-10, -1.342954e-08, -1.51469e-08, -1.084464e-08, -1.33893e-08, 
    -8.12912e-09, 7.3443e-08, -1.158213e-08, 2.445339e-07, -4.688576e-08, 
    3.673739e-08, 1.207906e-08, -6.319567e-11, 2.189773e-08, -1.445241e-07, 
    6.480703e-08, 3.498315e-09, -2.352587e-08, 8.568595e-09, 3.493625e-08, 
    -2.966857e-08, 6.037851e-09, -1.30528e-07, -4.376194e-08, -4.730978e-09, 
    -5.975198e-08, -1.284374e-07, 8.289859e-08, 1.974698e-08, -9.267154e-10, 
    -1.339629e-09, 1.015114e-07, 7.401934e-08, 8.168534e-08, 3.721212e-09, 
    -9.568453e-10, -3.842047e-10, 3.183288e-09, -1.675575e-08, -4.53305e-08, 
    -1.899099e-08, -6.515762e-08, 1.644702e-08, 7.539444e-08, -1.551206e-08, 
    -1.358567e-07, -8.929709e-08, 1.008459e-09, 8.977565e-09, -2.034799e-08, 
    -4.162473e-09, 9.419381e-10, -1.405667e-08, 2.180829e-09, -1.230298e-07, 
    5.665248e-08, 9.850382e-08, 2.360196e-09, -4.953904e-10, -1.132418e-08, 
    -9.157651e-08, -1.862394e-07, 2.788795e-09, 1.503888e-08, 3.901482e-08, 
    3.657249e-09, -5.723372e-09, 1.509648e-09, 1.148286e-07, -3.7034e-08, 
    3.002077e-08, -1.558144e-07, 9.489725e-09, -5.194863e-09, -1.452014e-08, 
    -1.696066e-08, -4.053192e-08, -1.830946e-08, 1.568218e-09, -3.323754e-08, 
    -2.409666e-08, -1.081031e-08, 3.138797e-08, 3.981307e-08, 3.29635e-10, 
    -7.490883e-09, -2.576712e-10, -2.862691e-09, -7.062397e-09, 
    -3.518039e-10, 9.178621e-10, -1.691802e-10, -3.74154e-10, 2.614087e-10, 
    2.930466e-08,
  1.457516e-08, -3.878426e-10, -1.336167e-08, -4.066686e-08, 3.361436e-09, 
    2.926794e-08, 9.426856e-09, -4.889955e-09, -9.554071e-09, -1.020356e-08, 
    -5.346635e-09, -1.374076e-09, -8.856262e-09, 2.727063e-09, -2.683697e-08, 
    3.321385e-08, -3.449684e-08, 4.37467e-10, 2.787338e-08, 8.208019e-09, 
    4.023815e-08, -5.597775e-08, 1.283013e-09, -3.309822e-09, 5.36204e-10, 
    9.072778e-10, -2.274766e-08, -9.527014e-09, -1.174629e-08, 4.103771e-08, 
    -1.258474e-08, -4.859822e-08, -6.005104e-08, 3.552939e-07, -7.251407e-08, 
    2.593043e-08, 1.356091e-08, -1.762714e-10, 2.447763e-08, -1.632315e-07, 
    3.165127e-08, 5.567415e-09, -1.341996e-07, 1.790379e-09, 3.073598e-08, 
    -1.328812e-08, 1.958711e-09, -1.391232e-07, -2.30864e-08, 8.837233e-10, 
    -6.051135e-08, -1.649574e-07, 8.012302e-08, 1.958573e-08, -4.98137e-09, 
    -2.597744e-10, 1.298666e-07, 7.79869e-08, 2.018281e-08, 1.441869e-08, 
    1.574165e-09, 1.985711e-09, 2.904301e-09, -1.534285e-08, -6.271087e-08, 
    -2.444364e-08, -5.924306e-08, 5.000408e-08, 4.998157e-08, -1.954066e-08, 
    -2.044591e-07, -3.510257e-08, 7.867641e-09, 9.524058e-09, -3.831474e-09, 
    1.227289e-08, 5.263459e-09, -1.487572e-08, 8.519692e-10, -1.428537e-07, 
    4.462669e-08, 1.786212e-07, 3.889056e-09, 5.377103e-09, -4.805258e-09, 
    -6.228623e-08, -2.644247e-07, 3.90429e-09, 1.678652e-08, 2.560489e-08, 
    -9.361543e-10, -1.993875e-09, 3.448122e-09, 1.463824e-07, -7.04361e-08, 
    6.517368e-08, -1.866577e-07, 4.674558e-08, -8.988366e-09, -1.271329e-08, 
    1.201645e-07, -3.759595e-08, -2.851259e-08, 2.616972e-09, -5.07502e-08, 
    -2.151666e-08, -3.976709e-09, 1.67235e-08, 6.350461e-08, 4.693163e-09, 
    -2.942613e-09, 5.03195e-09, -1.672902e-10, -2.666127e-09, 2.810907e-10, 
    5.252332e-11, -1.837321e-10, -1.051141e-09, 2.848566e-10, -2.970239e-09,
  1.680053e-08, -4.951062e-10, -3.448918e-09, -2.184572e-08, 1.154137e-08, 
    2.069271e-08, 8.293568e-09, 7.941026e-10, -3.829769e-09, -2.052047e-10, 
    3.718583e-09, 1.172225e-09, -8.222628e-09, -1.843034e-08, 2.043976e-09, 
    2.253569e-08, -5.233094e-08, 1.769638e-08, 5.730175e-08, 4.58806e-09, 
    6.002608e-08, -6.212815e-08, -1.126296e-09, -1.224066e-09, 6.156256e-09, 
    3.364528e-08, -2.290051e-08, 1.314436e-08, -1.676096e-08, 5.845698e-08, 
    -1.153433e-08, -5.928302e-08, -7.758592e-08, 1.519755e-07, -8.505447e-08, 
    -9.71329e-09, 6.471009e-09, -9.106316e-11, 4.122887e-08, -1.768451e-07, 
    1.790363e-09, 4.711069e-09, -2.658916e-07, -8.657963e-12, 2.112768e-08, 
    -3.185392e-09, 1.281023e-09, -1.665164e-07, -1.668743e-08, 1.679985e-08, 
    -5.468041e-08, -1.527152e-07, 8.921438e-08, 2.219129e-08, -8.959955e-09, 
    -1.61117e-09, 1.564759e-07, 5.649169e-08, -3.723162e-08, 1.869361e-08, 
    3.520313e-09, 1.778528e-08, -5.312245e-09, -4.680782e-09, -7.576143e-08, 
    -8.024813e-09, -3.833577e-08, 5.946083e-08, 1.879505e-08, -1.606361e-08, 
    -2.248938e-07, -4.405899e-08, 3.460912e-08, 1.435865e-10, 7.295967e-10, 
    4.641265e-09, 4.397663e-09, -8.900486e-09, -1.063154e-09, -8.105678e-08, 
    2.764205e-08, 2.001499e-07, 5.410016e-09, 5.111929e-09, -2.469164e-09, 
    -1.812634e-08, -4.432002e-08, 3.491323e-10, 1.486921e-08, 2.287777e-08, 
    3.483933e-09, -1.657487e-09, 4.993524e-09, 1.967029e-07, -6.890161e-08, 
    9.901746e-08, -1.743674e-07, 4.067181e-08, -1.106389e-08, -8.981329e-09, 
    4.268202e-08, -8.931266e-09, -2.118691e-08, 3.315307e-09, -6.72029e-08, 
    -1.601541e-08, 1.518799e-08, -8.432494e-09, 8.213885e-08, 1.197475e-08, 
    6.433538e-10, 1.42312e-08, 6.386131e-09, 7.289714e-09, 1.951662e-09, 
    -5.280298e-10, 4.218066e-10, -1.391307e-09, 3.174137e-10, -2.166269e-08,
  1.815897e-08, -2.237357e-09, 7.378276e-09, 4.416961e-09, 1.176454e-08, 
    1.839294e-08, 8.09905e-09, 2.501611e-08, 1.164494e-08, -3.718401e-08, 
    1.218041e-09, -5.979928e-11, -3.721129e-08, -3.954187e-08, 4.055391e-08, 
    -4.373556e-09, -5.966815e-08, 3.426635e-09, 8.522034e-08, -2.459637e-08, 
    3.913124e-08, -4.468802e-08, -1.826038e-09, -6.80302e-10, 7.070412e-09, 
    9.032487e-08, -1.810758e-08, 1.592389e-08, -1.979333e-08, 6.630466e-08, 
    1.058129e-08, -5.185871e-08, -7.17971e-08, 8.83756e-09, -9.229461e-08, 
    -2.159368e-08, -3.248556e-09, -1.556259e-09, 7.484664e-08, -1.843128e-07, 
    -4.485137e-08, -5.675247e-10, -2.619136e-07, 1.542253e-08, 1.772287e-08, 
    2.627257e-08, 1.507044e-08, -2.095241e-07, -1.60298e-08, 2.664214e-08, 
    -3.660438e-08, -1.205199e-07, 9.345124e-08, 3.196833e-08, -1.322542e-08, 
    1.300577e-10, 1.618666e-07, 2.99156e-08, -7.987899e-08, 1.151091e-08, 
    2.395382e-09, 3.597756e-08, -4.678668e-08, 2.879096e-08, -7.310305e-08, 
    2.980141e-08, -3.196647e-08, 1.836747e-08, -1.757735e-08, -6.440587e-09, 
    -1.525325e-07, -5.398033e-08, 2.226511e-07, -4.072035e-09, 9.781842e-10, 
    -3.183004e-09, 7.362843e-09, -2.817501e-09, -3.556863e-10, -3.875516e-08, 
    1.170451e-08, 1.648223e-07, 5.812922e-09, -3.14094e-09, -2.859224e-09, 
    -3.626383e-09, -7.802487e-08, -5.558604e-09, 1.472429e-08, 4.020933e-08, 
    8.218649e-09, 1.266606e-09, 2.456829e-09, 2.088036e-07, -6.166692e-08, 
    1.226858e-07, -1.294783e-07, 2.691581e-08, -1.349554e-08, -5.855918e-09, 
    -3.797732e-08, 1.619952e-08, -2.161819e-08, 2.859906e-09, -5.442075e-08, 
    4.509729e-08, 4.77371e-09, -8.131565e-09, 7.477934e-08, 1.385592e-08, 
    -4.151843e-10, 2.236629e-08, 1.502349e-08, 1.632293e-08, -1.503167e-09, 
    -1.094054e-09, 8.209895e-10, -1.44334e-09, 3.413874e-10, -1.112062e-08,
  1.610425e-08, -1.208861e-08, 1.79719e-08, 3.087342e-08, 6.346738e-09, 
    1.550171e-08, 1.451002e-08, 5.441535e-08, 2.539508e-08, -1.028163e-07, 
    -3.333508e-08, -1.899747e-08, -6.835859e-08, -5.77856e-08, 3.845133e-08, 
    -2.3704e-08, -7.882308e-08, -4.350227e-10, 1.096924e-07, -7.518128e-08, 
    5.094819e-09, -1.427844e-08, -6.277048e-09, -4.655476e-11, 3.582448e-08, 
    1.300085e-07, -6.52193e-09, 2.523558e-08, -1.718257e-08, 5.43734e-08, 
    8.192558e-09, -6.365161e-08, -5.703833e-08, -5.704266e-08, -9.268541e-08, 
    -1.824293e-08, -1.543889e-08, -1.377074e-09, 1.004506e-07, -1.785839e-07, 
    -9.982458e-08, -3.72637e-09, -1.194625e-07, 3.126316e-08, 9.22347e-09, 
    4.257862e-08, 1.558637e-07, -2.529516e-07, -1.718198e-08, 3.545112e-08, 
    -1.61053e-08, -1.246709e-07, 8.180967e-08, 3.907491e-08, -1.852302e-08, 
    2.103206e-11, 1.566643e-07, -9.460798e-08, -7.531341e-08, 1.070603e-08, 
    -1.284377e-09, -1.12571e-08, -1.053465e-07, 7.416878e-08, -5.878575e-08, 
    1.819052e-08, -3.001702e-08, -2.13675e-08, -4.374778e-08, 1.94683e-09, 
    -6.285347e-09, -2.610642e-08, 3.771145e-07, -5.67951e-09, 3.620516e-09, 
    -8.703239e-09, 1.439868e-08, 6.980883e-09, -7.970499e-10, -5.114867e-08, 
    -2.251284e-09, 1.203993e-07, 5.073844e-09, -1.877578e-08, 4.043443e-09, 
    -1.918465e-10, 1.196605e-08, -7.103097e-09, 3.136217e-08, 7.175214e-08, 
    6.692119e-09, 9.518558e-09, -8.947154e-11, 2.397263e-07, -5.531939e-08, 
    1.549294e-07, -6.964648e-08, -4.188036e-08, -2.123176e-08, -4.651804e-09, 
    7.071606e-09, 1.132509e-08, -1.979234e-08, 6.023448e-09, -6.476233e-08, 
    2.333053e-08, -5.935061e-08, 5.478284e-09, 4.550935e-08, 7.130382e-09, 
    -7.120832e-09, 2.120163e-08, 1.243671e-08, 1.225027e-08, -1.116047e-08, 
    -7.627364e-10, 2.829694e-09, -1.481034e-09, 3.846878e-10, -9.535199e-09,
  1.247963e-08, -3.424793e-08, 7.216386e-09, 3.448622e-08, -3.819423e-09, 
    3.455625e-09, 1.522812e-08, 4.710569e-08, 3.624336e-08, -7.516746e-08, 
    -7.996164e-08, -4.587264e-09, -3.234413e-08, -5.010202e-08, 7.217295e-09, 
    -1.722158e-08, -5.818838e-08, -7.838025e-09, 2.148431e-08, -1.729222e-07, 
    -8.325287e-08, 5.181846e-09, -1.998592e-08, 1.690228e-08, 4.387744e-08, 
    7.690255e-08, 1.287867e-08, 2.975776e-08, -1.66342e-08, 9.021505e-09, 
    -1.712465e-08, -8.683537e-08, -6.138521e-08, -1.370659e-07, 
    -7.735525e-08, -1.568992e-08, -2.016473e-08, -1.919233e-09, 1.130757e-07, 
    -1.7077e-07, -1.462213e-07, -8.508778e-09, 1.629479e-08, 3.211142e-08, 
    -2.049319e-09, 1.669241e-08, 5.843663e-08, -3.12055e-07, -3.69485e-08, 
    3.5089e-08, -6.52463e-09, -1.577348e-07, 5.202178e-08, 4.107142e-08, 
    -2.562868e-08, 3.072955e-10, 1.451217e-07, -1.224503e-07, -4.293268e-08, 
    3.638544e-08, -3.393325e-09, 1.676628e-07, -1.201574e-07, 1.218151e-07, 
    -3.490977e-08, 2.57146e-08, -3.037076e-08, -3.943023e-08, -7.114977e-08, 
    1.092553e-08, 4.63483e-08, 7.119752e-09, 8.512711e-08, -6.723894e-09, 
    1.409498e-08, -2.015918e-08, 5.577817e-09, 1.194553e-08, -4.934361e-09, 
    -9.565542e-08, -1.709975e-08, 7.574991e-08, 3.570221e-09, -2.642992e-09, 
    2.022716e-09, 3.520404e-08, 6.861455e-09, -1.209128e-08, 5.302646e-08, 
    8.781785e-08, 1.226203e-08, 1.438021e-08, -4.236426e-09, 2.842966e-07, 
    -7.943754e-09, 2.046961e-07, -2.317766e-08, -3.994342e-08, -3.47793e-08, 
    -2.235356e-09, 3.209811e-08, -1.566895e-08, -2.710043e-08, 1.405394e-08, 
    -8.293227e-08, -2.26903e-08, -7.210429e-08, 4.576123e-09, 5.708443e-09, 
    -2.328079e-09, -2.445313e-08, 8.600864e-09, -5.026095e-09, 2.028946e-08, 
    -1.172134e-08, -3.401283e-10, 2.87551e-09, -1.305914e-09, 4.862386e-10, 
    1.305727e-07,
  7.589506e-09, -6.055166e-08, -3.103446e-08, 4.936965e-09, 6.170922e-10, 
    -5.666152e-09, 1.217586e-08, 3.216519e-08, 4.362619e-08, -3.50808e-08, 
    -6.873029e-08, 3.478683e-07, -2.243723e-08, -3.796094e-08, -3.919399e-08, 
    -2.048864e-09, -4.230695e-08, -1.604576e-09, 2.288448e-08, -1.052256e-07, 
    -2.443721e-07, 5.078755e-08, 1.382466e-07, 5.667732e-07, 6.964001e-08, 
    6.46537e-08, 3.536707e-08, 2.489173e-08, 1.214721e-08, -6.82121e-10, 
    -5.180027e-09, -1.19695e-07, -6.039841e-08, -1.932613e-07, -7.038216e-08, 
    -4.028652e-08, -1.676749e-08, -3.157595e-09, 1.129165e-07, -1.464837e-07, 
    -1.376277e-07, -5.620677e-09, 1.199487e-08, 4.2125e-08, -1.647823e-08, 
    -2.63924e-08, 4.896833e-09, -3.621231e-07, -2.968495e-08, 3.183284e-08, 
    3.304245e-08, -2.491593e-07, 2.24597e-08, 4.43677e-08, -3.236539e-08, 
    5.337597e-10, 1.398539e-07, -4.866213e-08, -1.635847e-08, 7.201535e-08, 
    -2.771458e-09, -5.618153e-08, -9.610562e-08, 1.483603e-07, -2.867336e-08, 
    2.715592e-08, -3.661376e-08, -3.014088e-08, -7.666381e-08, 1.97947e-08, 
    8.023085e-08, 4.849358e-08, 4.207413e-08, -9.000587e-09, 4.689955e-08, 
    -1.674334e-08, -2.504066e-09, 1.452855e-08, -1.099562e-08, -1.302185e-07, 
    -3.733692e-08, 3.514815e-08, 2.499974e-09, -1.59223e-08, -1.416856e-08, 
    1.007329e-07, -9.935729e-08, -2.425327e-08, 3.983028e-08, 8.511643e-08, 
    3.111586e-08, -1.573561e-09, -1.45352e-08, 2.836516e-07, -4.752337e-09, 
    2.022731e-07, -4.194999e-09, 5.096467e-08, -4.196795e-08, 1.609892e-08, 
    5.084962e-08, -6.288739e-08, -3.922686e-08, 2.16961e-08, -8.128836e-08, 
    -4.885646e-08, -2.996717e-08, 8.08086e-10, -2.790239e-08, -1.838816e-08, 
    -4.556955e-08, 1.439957e-09, -8.340066e-09, 4.302842e-08, -5.627044e-09, 
    -8.774805e-10, 9.76911e-10, -1.219775e-09, 5.860699e-10, 1.021874e-07,
  6.204289e-09, -7.300793e-08, -9.377601e-08, -3.601377e-08, 1.448637e-08, 
    5.960771e-09, 1.282746e-08, 3.066901e-08, 5.42388e-08, -1.591826e-08, 
    -4.79809e-08, -1.881659e-08, 4.912806e-09, -3.440624e-08, 5.494428e-09, 
    3.652837e-09, -3.892843e-08, 1.643514e-09, 8.253005e-08, 5.500794e-09, 
    -2.438383e-07, 2.898966e-07, -2.194594e-08, -7.957743e-08, 1.76026e-07, 
    4.086377e-08, 3.068106e-08, 2.537257e-08, 2.734618e-08, 1.841789e-08, 
    3.339932e-08, -7.332875e-08, -4.793066e-08, -1.777822e-07, -4.328928e-08, 
    -6.357965e-08, -2.543732e-09, -3.056158e-09, 1.076291e-07, -1.160891e-07, 
    -3.607411e-08, 2.614785e-07, -1.017423e-07, 5.209578e-08, -1.214477e-08, 
    -5.17087e-08, -1.37299e-08, -4.01913e-07, -3.279839e-08, 2.585482e-08, 
    3.440954e-08, -6.679448e-08, -1.028214e-08, 5.451606e-08, -3.775858e-08, 
    3.507807e-10, 1.129194e-07, -1.591965e-08, 1.28781e-09, 1.282549e-07, 
    -1.241062e-09, -4.552777e-08, -5.880798e-08, 1.215648e-07, -4.978685e-08, 
    2.86779e-08, -4.039913e-08, -1.705968e-08, -5.973658e-08, 1.798998e-08, 
    9.149511e-08, 9.815784e-08, 7.412285e-08, -3.81238e-08, 1.235256e-07, 
    -1.116797e-08, -4.296169e-09, 1.240221e-08, -1.517489e-08, -9.758247e-08, 
    -5.249223e-08, 1.229403e-08, 3.076195e-09, -1.234696e-09, -1.32805e-08, 
    2.89121e-08, -9.90147e-08, -1.23635e-08, 1.473515e-08, 6.189561e-08, 
    5.821147e-08, -2.946619e-08, -1.647714e-08, 2.345166e-07, -1.686755e-08, 
    1.740709e-07, 6.801569e-08, -4.7573e-08, -4.347686e-08, 1.691877e-08, 
    7.021976e-08, -1.075779e-07, -5.015495e-08, 2.089844e-08, 4.779616e-08, 
    -5.636576e-08, 2.748033e-08, -2.15465e-09, -4.823943e-08, -3.610177e-08, 
    -4.062514e-08, -4.066635e-09, 1.74208e-09, 6.085378e-08, -3.184425e-09, 
    -1.44604e-09, 1.376321e-09, -9.9039e-10, 6.634622e-10, 1.002597e-07,
  4.838682e-09, -5.813041e-08, -1.108329e-07, -6.274655e-08, 1.482084e-08, 
    2.713494e-08, 2.574797e-08, 6.416093e-08, 4.359293e-08, -1.034851e-08, 
    -1.1753e-08, -9.676575e-08, -9.243706e-09, -4.206009e-08, -3.875749e-08, 
    6.17141e-09, -3.318043e-08, 2.165399e-08, 5.128078e-08, 7.454759e-08, 
    -4.335612e-08, 1.250595e-08, -3.459155e-08, -1.003951e-07, 4.014241e-07, 
    -8.410649e-08, 3.845724e-08, 3.045551e-08, 1.351617e-08, 2.518908e-08, 
    6.197678e-08, -2.604571e-08, -1.850759e-08, -1.087206e-07, -1.581213e-09, 
    -5.384101e-08, 1.021657e-08, -2.904358e-09, 9.604531e-08, -1.035039e-07, 
    -4.839586e-08, 1.325651e-08, -1.479922e-07, 4.904666e-08, 5.56696e-09, 
    -4.281816e-08, -2.146118e-08, -4.009185e-07, -2.391445e-08, 1.818655e-08, 
    3.526864e-08, -6.235251e-08, -3.078697e-08, 6.361669e-08, -4.365072e-08, 
    -1.197293e-09, 8.937849e-08, 4.527248e-09, 4.283436e-09, 2.370999e-07, 
    2.386457e-09, 2.285509e-08, 1.902725e-08, 9.110412e-08, -3.192574e-08, 
    3.700092e-08, -4.314558e-08, -1.576211e-09, -4.617465e-08, 1.514121e-08, 
    8.567866e-08, 1.159048e-07, 6.733961e-08, -5.76286e-08, 9.889046e-08, 
    -6.722587e-09, 1.385806e-08, 1.405419e-08, -1.796483e-08, -3.582642e-08, 
    -6.077875e-08, 1.74761e-08, 8.476434e-09, 5.856504e-08, -4.911328e-09, 
    9.194758e-08, -9.320053e-08, 4.596984e-09, 3.399285e-08, 2.937367e-08, 
    -1.611973e-07, -3.776537e-08, -3.318462e-09, 1.894268e-07, -2.690132e-08, 
    2.10884e-07, 9.071472e-08, -4.996019e-08, -3.626093e-08, -1.933702e-10, 
    1.920727e-07, -1.055625e-07, -5.978677e-08, 1.161386e-08, 5.027545e-08, 
    -1.530208e-08, 5.014675e-08, -9.523376e-09, -5.789462e-08, -4.57315e-08, 
    -2.688972e-08, -1.441532e-08, 2.413543e-08, 5.839155e-08, -1.269257e-09, 
    -1.666706e-09, 2.388845e-10, -8.06665e-10, 6.786252e-10, -4.879467e-08,
  7.185008e-10, -1.72779e-08, -6.026903e-08, -4.204549e-08, 2.944262e-09, 
    6.852474e-08, 7.113204e-08, 1.360374e-07, 1.243052e-08, -1.711305e-08, 
    1.102771e-07, -1.152778e-07, -2.201818e-08, 3.135915e-08, -2.035613e-07, 
    1.148759e-09, -2.684394e-08, 8.589382e-09, 8.503315e-08, 1.179001e-07, 
    -1.064109e-10, -9.198629e-09, 3.376567e-08, -3.315199e-08, -1.709805e-08, 
    -1.443066e-07, 5.883271e-08, 3.15938e-08, -1.289072e-08, 2.964816e-08, 
    9.445603e-08, -1.548665e-08, -2.501861e-08, -4.419735e-08, 1.754529e-08, 
    -2.150068e-08, 1.696369e-08, -2.74278e-09, 7.322546e-08, -1.017352e-07, 
    -5.780579e-08, -1.16479e-08, -1.213645e-07, 4.248407e-08, -1.75653e-08, 
    -4.091021e-08, -1.329737e-07, -2.963852e-07, -2.07599e-08, 9.445685e-09, 
    3.55671e-08, -6.196933e-08, -4.138785e-08, 6.667428e-08, -5.247146e-08, 
    -6.932282e-09, 7.183849e-08, 1.085293e-08, 6.878108e-08, 3.428511e-07, 
    3.437435e-09, -1.094088e-07, 9.294808e-08, 6.352474e-08, -9.874839e-09, 
    2.670072e-08, -2.162756e-08, -8.27481e-09, -4.510252e-08, 4.066806e-09, 
    7.463632e-08, 9.45488e-08, 2.603497e-08, -4.606272e-08, -5.667132e-08, 
    -3.510877e-09, 9.33349e-09, 1.311736e-08, -2.376717e-08, -7.407243e-08, 
    -7.02795e-08, 2.170678e-08, -2.261004e-09, 2.448594e-07, 7.428525e-09, 
    9.789119e-09, -1.297828e-07, 8.633378e-09, 5.686788e-08, -1.198828e-09, 
    3.874766e-08, -3.984988e-08, -2.686704e-09, 1.695885e-07, -1.559761e-08, 
    2.335166e-07, 7.054773e-08, -5.515199e-08, -6.75891e-09, -2.904653e-09, 
    1.789317e-08, -1.104966e-07, -6.647807e-08, 3.640849e-09, 2.577485e-08, 
    1.572243e-08, 3.352011e-08, -2.025399e-08, -6.663777e-08, -4.962362e-08, 
    -2.257548e-08, -1.401054e-08, 2.925822e-08, 2.282377e-08, -1.321519e-08, 
    -5.406942e-11, 2.775096e-09, -3.418158e-09, 7.281358e-10, -4.194044e-08,
  -8.639063e-10, 3.166076e-08, -4.126491e-09, -2.13937e-08, -4.51347e-08, 
    1.818536e-07, 1.650168e-07, 3.422537e-07, -1.252135e-08, 3.241269e-08, 
    -7.226538e-08, -2.485115e-08, 1.899886e-07, -6.11293e-08, -1.670861e-07, 
    -4.001231e-09, 4.12129e-09, 6.673167e-08, 5.704828e-08, 1.589032e-07, 
    -4.932156e-08, 3.785772e-11, 2.711602e-08, -4.141725e-09, 1.902879e-08, 
    -7.134247e-08, 5.66987e-08, 2.88079e-08, -4.084143e-08, 1.380465e-08, 
    1.476373e-07, -3.853359e-08, 8.534369e-08, -7.566655e-09, 2.138165e-08, 
    -3.302455e-08, 2.75754e-08, -2.093856e-09, 4.315245e-08, -1.095163e-07, 
    -5.764753e-08, -2.463855e-08, -5.454427e-08, 3.914544e-08, -1.481737e-08, 
    -4.609058e-08, -1.456993e-07, -2.430725e-07, -1.918254e-08, 2.318146e-09, 
    3.621952e-08, -2.369109e-08, -3.959251e-08, 6.63382e-08, -4.425874e-08, 
    -3.432319e-09, 5.317327e-08, -1.521723e-08, 3.117993e-07, 9.667502e-08, 
    1.690063e-07, -1.466693e-07, 3.381126e-08, 2.949084e-08, 1.532187e-08, 
    2.86833e-08, -2.405216e-08, -2.436911e-08, 6.378627e-09, -4.62785e-09, 
    6.272728e-08, 5.454433e-08, -2.962122e-08, 5.191737e-09, -6.357084e-08, 
    1.385274e-09, 1.419693e-09, 1.772486e-08, -1.773159e-08, -2.893523e-08, 
    -8.906807e-08, 4.454161e-08, -9.690893e-09, 1.098093e-07, 1.72671e-08, 
    3.794196e-08, -1.019038e-07, 2.239972e-09, 7.440508e-08, -1.600552e-08, 
    2.972558e-08, -2.964173e-08, -6.549442e-09, 1.551057e-07, 4.527806e-09, 
    2.568179e-07, 4.31857e-08, -6.805647e-08, 1.619549e-08, -2.642553e-08, 
    -7.561846e-08, 1.341624e-08, -7.100763e-08, -1.384237e-09, -1.234378e-08, 
    2.101444e-08, 2.798981e-08, -3.03188e-08, -7.378401e-08, -5.213553e-08, 
    -1.956585e-08, -1.137676e-08, 7.302901e-09, -1.612614e-08, -5.420475e-09, 
    1.544913e-09, 2.422524e-09, -2.093053e-09, -5.934027e-10, -6.400012e-08,
  7.811082e-09, 8.028394e-08, -1.636056e-08, -1.639756e-07, 5.329741e-08, 
    4.204693e-07, 2.411286e-08, -5.572758e-08, 1.440097e-07, 1.598698e-08, 
    -8.485006e-08, 5.832476e-09, -3.700882e-08, -9.314601e-08, -2.405602e-08, 
    -7.090444e-09, 3.675495e-08, 8.810514e-08, 7.698119e-08, 7.8786e-08, 
    4.536673e-09, 1.908813e-08, 1.268799e-07, 1.226942e-08, 8.76463e-08, 
    1.838873e-08, 6.748417e-08, 2.250806e-08, -6.298035e-08, -4.589879e-09, 
    1.585944e-07, 9.361315e-09, 1.946636e-07, 1.643343e-09, 3.489856e-08, 
    -4.121819e-08, 4.090766e-08, -1.308905e-09, 1.642036e-08, -1.304277e-07, 
    -5.319059e-08, -9.172766e-08, -7.247883e-08, 3.850543e-08, -2.631293e-08, 
    -8.861036e-08, -9.759208e-08, -2.364069e-07, -2.35879e-08, -1.716955e-10, 
    3.600923e-08, -9.993857e-08, -2.177169e-08, 6.236525e-08, -2.972654e-08, 
    -6.093615e-11, 3.951038e-08, -1.797867e-09, 4.238983e-07, 6.914516e-08, 
    -1.997881e-07, -1.127984e-07, 2.321951e-08, 2.247368e-08, 4.988726e-08, 
    2.887475e-08, -3.655828e-09, -3.570733e-08, 2.37593e-08, -1.227875e-08, 
    3.345906e-08, 1.939611e-09, -9.066241e-08, -1.405067e-08, -4.032859e-08, 
    5.853167e-09, 2.866756e-09, 1.817165e-08, -2.427871e-08, 1.985165e-08, 
    -1.114161e-07, -1.768294e-08, -1.481794e-08, 3.53017e-08, 5.63449e-08, 
    8.847678e-09, -6.589778e-08, -7.302901e-09, 6.671138e-08, -1.526428e-08, 
    1.295972e-07, -1.569149e-08, -5.082086e-09, 1.277915e-07, -1.543833e-08, 
    2.671679e-07, 2.144e-08, 3.759624e-10, 1.626961e-08, -1.933153e-09, 
    -1.840669e-08, -5.584734e-08, -7.054956e-08, -2.334389e-09, 
    -1.398428e-08, -1.587625e-08, 3.243179e-08, -3.919865e-08, -7.957067e-08, 
    -5.418326e-08, -1.838941e-08, -1.056799e-08, -3.169021e-09, 
    -1.043088e-08, 2.053525e-09, 3.154264e-09, 1.956494e-09, -2.314827e-09, 
    -4.194618e-10, -2.54571e-08,
  1.193501e-08, 1.197653e-07, -6.070642e-07, -5.99439e-07, -8.132264e-08, 
    1.285917e-07, 5.79206e-09, -1.355062e-08, 1.412224e-08, -2.478401e-08, 
    -3.243025e-08, 8.445892e-08, -2.493329e-08, -2.013581e-08, 3.150092e-09, 
    -2.349614e-08, 4.972929e-08, 6.962574e-08, 7.055415e-08, 8.838299e-09, 
    7.243392e-08, 3.008603e-08, 1.41676e-08, -6.456713e-08, -1.795598e-08, 
    5.016892e-08, 5.43186e-08, 2.0198e-08, -6.861097e-08, -2.811873e-09, 
    1.168984e-07, -1.535096e-08, 7.637055e-08, 4.269509e-10, 3.70531e-08, 
    -2.314647e-08, 5.085145e-08, -1.290559e-09, -4.237847e-09, -1.480617e-07, 
    -1.444915e-08, -9.211789e-08, -9.329818e-08, 4.684824e-08, -1.882137e-08, 
    -8.966566e-08, -7.238413e-08, -1.465932e-07, -1.499785e-08, 4.855991e-10, 
    3.573135e-08, -9.612637e-08, 3.621289e-09, 5.823512e-08, -2.938762e-08, 
    -7.143512e-10, 2.761254e-08, 1.357532e-08, 9.539148e-08, 1.487502e-07, 
    -1.613817e-07, -8.728222e-08, 1.351655e-07, 1.105115e-08, 8.749357e-08, 
    2.277187e-08, 5.740668e-08, -3.618521e-08, 9.32954e-09, -2.176529e-08, 
    5.898642e-10, -2.647454e-08, -1.306126e-07, -5.735791e-08, -3.285408e-10, 
    5.105392e-09, 4.844864e-09, 2.104605e-08, 3.219284e-09, -1.407119e-08, 
    -1.212103e-07, -4.7083e-09, -2.355006e-08, -1.042532e-07, 9.575245e-08, 
    -5.050839e-08, -3.232515e-09, -2.108624e-08, 5.371135e-08, -2.31496e-08, 
    4.613906e-08, -2.433677e-08, 9.332837e-10, 7.489855e-08, 1.727415e-09, 
    2.671175e-07, 1.519005e-08, 1.546181e-08, 3.20087e-08, 4.922243e-09, 
    1.093917e-07, -6.960367e-08, -7.546137e-08, -4.036877e-09, -2.540065e-08, 
    -5.214946e-08, 4.614895e-08, -4.802399e-08, -8.475098e-08, -5.589192e-08, 
    -1.789937e-08, -9.191638e-09, -3.358252e-09, 2.508216e-09, 2.964555e-09, 
    3.677053e-09, 2.464105e-09, -2.594792e-09, -2.427143e-10, -1.310906e-07,
  5.023736e-08, 3.627764e-08, -1.100156e-06, -1.464423e-07, -4.567181e-08, 
    2.020153e-08, -2.191825e-09, -1.177756e-08, -6.250144e-08, -1.799407e-08, 
    -3.365273e-08, 9.112892e-08, -2.555197e-08, 1.899178e-08, 3.610296e-09, 
    -3.538164e-08, 5.514842e-08, 3.27438e-08, 1.940454e-08, -7.665847e-09, 
    2.238352e-07, -1.963662e-08, 7.547959e-08, -1.197748e-09, -5.807863e-09, 
    6.424403e-08, 1.413326e-08, 1.29366e-08, -5.712417e-08, 4.198625e-09, 
    6.582439e-08, 5.410544e-08, -7.77078e-09, -7.946545e-08, 2.069868e-08, 
    2.033027e-07, 5.924219e-08, -1.634703e-09, -1.596931e-08, -1.544684e-07, 
    5.591995e-08, 2.086114e-08, -3.851392e-08, 4.919672e-08, -2.785686e-08, 
    -1.209058e-07, -5.644847e-08, -9.003628e-08, -2.457367e-08, 2.122249e-09, 
    3.532756e-08, 5.748569e-08, 1.917381e-08, 4.694672e-08, -2.504898e-08, 
    -1.190926e-09, 2.9668e-08, 1.567412e-08, -7.65753e-08, 1.955291e-08, 
    -3.751251e-08, -3.112513e-08, -9.638939e-10, -1.564887e-08, 9.413029e-08, 
    1.175687e-08, 8.125056e-08, -2.200892e-08, 5.438511e-08, -3.337158e-08, 
    -7.070582e-09, -5.619938e-09, -1.334419e-07, -6.209171e-08, 2.116558e-09, 
    9.442886e-09, 2.239889e-08, 9.180297e-09, 2.307972e-08, 5.813951e-08, 
    -1.121025e-07, 9.533551e-09, -3.281417e-08, -3.432637e-07, 7.928321e-08, 
    -3.530164e-08, 9.938645e-08, -5.84302e-08, 2.000698e-08, -1.519351e-08, 
    -2.2395e-08, -3.146475e-08, 9.854261e-09, 5.737324e-08, 1.30953e-08, 
    2.683435e-07, 8.059773e-09, 2.791415e-08, 4.867496e-08, 2.221008e-08, 
    1.575415e-07, -4.794373e-09, -9.84865e-08, -5.294247e-09, -4.57872e-08, 
    -2.578059e-08, 6.681222e-08, -5.680425e-08, -8.935234e-08, -5.850205e-08, 
    -1.73755e-08, -9.362395e-09, -4.708284e-09, 5.002505e-09, 2.509807e-09, 
    5.040124e-09, 3.021341e-09, -2.638515e-09, 2.357154e-10, -1.401312e-07,
  -1.38229e-08, -5.149209e-07, -1.916735e-07, 9.216473e-08, -4.070995e-08, 
    -1.41037e-07, 1.421262e-08, 1.283132e-08, 9.956182e-09, -2.301528e-08, 
    -3.451947e-08, 8.188664e-08, 1.444818e-08, -1.107827e-08, 5.106074e-09, 
    -1.552666e-08, 6.080376e-08, 3.142031e-08, -3.790947e-08, -6.324871e-08, 
    2.488861e-08, -1.616132e-08, 7.269222e-08, 7.669883e-10, -1.672839e-08, 
    1.459458e-07, -7.082525e-08, 1.084965e-08, -3.830024e-08, -9.406165e-09, 
    -6.895959e-09, 7.546561e-08, -4.520365e-08, -2.474468e-08, -4.461896e-08, 
    1.514687e-07, 6.858929e-08, -1.112085e-09, -1.256745e-08, -1.232834e-07, 
    1.276756e-07, 3.436713e-08, 5.459194e-08, 2.849926e-08, -2.291785e-08, 
    -7.537511e-08, -5.377291e-08, -6.731531e-08, -3.586819e-08, 3.746699e-09, 
    3.478358e-08, 3.770672e-07, 2.228718e-08, 3.360459e-08, -2.366384e-08, 
    -4.176286e-09, 3.426106e-08, 5.058027e-08, -9.244909e-08, -8.275649e-09, 
    -1.073869e-08, 2.512701e-08, 1.503525e-08, 1.093773e-08, 7.181785e-08, 
    3.333241e-09, 9.608613e-08, -1.122714e-09, 1.706127e-08, -2.971564e-08, 
    -5.155982e-09, -5.520332e-08, -1.884592e-08, -1.705968e-08, 
    -6.709939e-09, 1.132383e-08, 6.556432e-08, 1.831893e-08, -2.407029e-09, 
    5.635349e-08, -9.098358e-08, 2.886266e-08, -5.397544e-08, -4.705475e-07, 
    2.761686e-08, 5.106148e-08, 5.427859e-08, -1.095105e-07, -1.143824e-08, 
    -7.568076e-09, -1.503793e-09, -2.720889e-08, 9.723777e-09, 4.923741e-08, 
    4.363215e-07, 2.667713e-07, 1.053003e-09, -1.453208e-08, -9.852045e-09, 
    5.832006e-08, 1.018549e-08, 3.310497e-09, 8.830256e-09, -3.807699e-09, 
    -2.698414e-09, 2.819945e-09, 8.273304e-08, -6.583156e-08, -9.503054e-08, 
    -6.181284e-08, -1.699385e-08, -9.655139e-09, -4.944752e-09, 5.214872e-09, 
    1.933643e-09, 5.051902e-09, 3.086569e-09, -1.790902e-09, 2.321983e-10, 
    -3.167764e-08,
  -4.454648e-09, -5.097724e-07, 6.019758e-08, 1.155644e-07, -8.221087e-08, 
    -1.415377e-07, 1.190659e-08, -4.334311e-10, 2.473541e-09, -1.76862e-08, 
    1.695088e-08, 7.253192e-08, -6.423022e-09, -1.256916e-08, -2.209902e-09, 
    5.226945e-09, 5.693488e-08, 3.9898e-08, 1.139232e-08, -2.173422e-07, 
    -6.027108e-10, -1.41336e-08, 7.360433e-08, 2.999684e-09, -2.660278e-08, 
    4.172028e-08, -9.570778e-08, 6.011135e-09, -3.27405e-08, -4.703355e-08, 
    -4.615134e-08, 7.63369e-08, 2.146675e-08, -3.03782e-08, 2.35479e-08, 
    1.451758e-07, 7.742916e-08, -8.223822e-11, 9.130929e-09, -1.006725e-07, 
    1.407333e-07, 3.897986e-08, 2.107643e-08, 2.53657e-08, -7.533515e-09, 
    -7.06562e-08, -5.492382e-08, -5.44814e-08, -3.366825e-08, 4.663569e-09, 
    3.409438e-08, -4.562679e-08, 2.255166e-08, 2.888113e-08, -2.280691e-08, 
    -4.110291e-09, 1.762038e-08, 8.335075e-08, -1.486133e-07, 1.901796e-09, 
    -9.063285e-09, 3.288352e-08, 1.682014e-08, 6.224957e-09, 4.917196e-08, 
    -1.351174e-08, 5.875262e-08, 1.043173e-08, 1.042855e-08, -3.102951e-08, 
    -8.728705e-09, -1.172127e-07, 2.011051e-07, -1.265283e-08, -1.277812e-08, 
    -6.326673e-11, -2.159142e-08, 1.578826e-08, -8.087349e-09, 2.219122e-07, 
    -7.139874e-08, 1.736771e-08, -7.392043e-08, -9.250414e-09, 2.118156e-09, 
    1.653834e-07, 4.764348e-08, -7.173941e-08, -2.704857e-08, -1.724231e-09, 
    1.293466e-08, -1.805623e-08, -1.268461e-09, 5.26927e-08, 3.866396e-07, 
    2.721457e-07, 6.513496e-09, -1.806231e-07, -8.016116e-09, 1.061163e-08, 
    -1.153912e-07, 6.375835e-09, 5.642086e-09, -3.76027e-09, -4.232828e-08, 
    -1.392988e-08, 9.552338e-08, -8.140086e-08, -1.066084e-07, -6.541023e-08, 
    -1.684788e-08, -9.926282e-09, -4.177252e-09, 5.155186e-09, 1.754245e-09, 
    3.82513e-09, 4.082779e-09, -1.241705e-09, -1.999751e-10, 3.156896e-08,
  -3.930671e-08, -8.35343e-08, 6.94759e-08, -3.717781e-08, -1.446068e-08, 
    -8.26837e-08, 4.797187e-09, 1.380442e-09, 7.720757e-09, 1.178768e-08, 
    -7.010783e-09, 1.108043e-07, -4.796505e-09, -1.324094e-08, -3.466255e-09, 
    1.317582e-08, 6.808999e-08, 2.32456e-08, 2.042512e-08, -1.018064e-07, 
    -1.019356e-08, -1.259917e-08, 7.368266e-08, 4.06402e-09, -2.667747e-08, 
    -4.823903e-09, -4.733084e-08, 7.949723e-09, -4.918439e-08, -7.23191e-08, 
    -1.255175e-07, 1.951188e-07, 4.944997e-08, 1.452958e-08, 3.156862e-08, 
    9.235163e-08, 7.939667e-08, 6.530456e-10, 4.760187e-08, -9.750801e-08, 
    1.68171e-07, 4.082273e-08, -4.961839e-08, 4.412158e-09, -4.53673e-09, 
    -7.655439e-08, -5.777048e-08, -5.224021e-08, -3.313668e-08, 5.689692e-09, 
    3.325241e-08, -6.127874e-08, 1.871355e-08, 2.333869e-08, -2.228404e-08, 
    -2.609909e-09, -1.978373e-08, 9.498076e-08, -1.877967e-07, -7.984156e-09, 
    -1.04356e-08, 3.977385e-08, 1.72252e-08, -5.078948e-09, 4.874356e-08, 
    -3.001145e-08, 1.761367e-08, 1.150721e-08, -2.541071e-09, -5.796136e-08, 
    1.51818e-08, -1.229456e-07, -3.689735e-08, -2.968761e-09, -1.815231e-08, 
    8.128552e-09, -1.256083e-09, 1.457374e-08, -1.260522e-08, -4.439931e-08, 
    -5.919719e-08, 1.457097e-08, -1.064674e-07, 4.913005e-08, 2.932723e-09, 
    1.773805e-08, 6.537351e-08, 9.883081e-09, -3.785065e-08, -1.368392e-09, 
    1.405425e-08, -1.367088e-08, -4.107875e-09, 5.349222e-08, 2.905477e-08, 
    2.843685e-07, 2.413833e-09, -3.549965e-07, -5.504097e-08, -1.147508e-08, 
    -8.704075e-08, 7.417512e-09, 3.365024e-09, -5.526694e-09, -1.957628e-07, 
    2.423292e-09, 1.084076e-07, -6.700492e-08, -7.686828e-08, -7.10865e-08, 
    -1.673646e-08, -1.026552e-08, -2.881904e-09, 5.005006e-09, 2.747754e-09, 
    4.529647e-09, 4.365802e-09, -2.324285e-09, 2.610605e-10, 4.441728e-08,
  -1.148099e-07, -6.344618e-08, 2.81795e-08, -6.309295e-08, 1.02587e-08, 
    -4.998952e-08, 4.534229e-09, 1.558135e-09, 8.055224e-09, 1.365055e-08, 
    -1.977298e-09, 8.262526e-08, -1.458545e-09, -1.301754e-08, 4.008655e-09, 
    8.232302e-09, 7.38162e-08, -2.569607e-09, 2.33875e-08, -7.848388e-08, 
    -1.44525e-08, -1.309417e-08, 7.494231e-08, 4.655988e-09, -2.447877e-08, 
    -2.426003e-08, 2.627581e-08, 4.220436e-08, -8.220383e-08, 3.242002e-08, 
    -1.129835e-07, 6.506906e-08, -8.121509e-08, 6.171018e-08, 3.236113e-08, 
    5.330691e-08, 7.449702e-08, 7.311343e-10, 4.296277e-08, -8.474213e-08, 
    1.675512e-07, 4.139548e-08, -8.366806e-08, 3.691179e-08, 3.701717e-08, 
    -6.737054e-08, -5.847755e-08, -5.534358e-08, -1.710138e-08, 6.542962e-09, 
    3.233728e-08, -6.579461e-08, 1.331622e-08, 1.966931e-08, -2.195561e-08, 
    -1.867988e-09, -5.859073e-08, 1.041882e-07, -2.188631e-07, -5.337782e-09, 
    -1.376122e-09, 4.323289e-08, 1.680434e-08, -3.108823e-09, 5.568906e-08, 
    -8.105638e-08, -1.279147e-09, -1.705587e-09, -3.475571e-08, 
    -5.284761e-08, 6.155352e-08, -1.247051e-07, -6.924614e-08, 9.013661e-10, 
    -2.186084e-08, 6.275229e-09, 1.394e-09, 4.909793e-09, -1.609218e-08, 
    -4.93863e-08, -3.55866e-08, 2.059219e-08, -1.097909e-07, 6.240424e-08, 
    3.17101e-09, 4.242281e-09, 1.287597e-07, 4.101764e-09, -4.604505e-08, 
    -4.575384e-09, 1.39309e-08, -5.084269e-09, -5.441848e-09, 4.976574e-08, 
    -6.630938e-08, 2.995833e-07, -1.421973e-08, -9.340403e-08, -6.086594e-08, 
    2.989395e-10, -5.905861e-09, 8.748891e-09, 1.79962e-09, -6.059999e-09, 
    -2.840977e-09, 3.531835e-08, 1.157683e-07, -2.1478e-08, -4.776524e-08, 
    -5.787064e-08, -1.568202e-08, -1.038023e-08, -1.979004e-09, 4.84971e-09, 
    1.33997e-09, 2.803858e-09, 5.724559e-10, -1.21598e-09, 5.24885e-10, 
    5.008593e-08,
  -8.023841e-08, -5.825206e-08, 2.746373e-08, -6.388046e-08, 1.379357e-08, 
    -2.630401e-08, 5.008985e-09, 2.900322e-09, 7.654023e-09, 9.214261e-09, 
    -2.444324e-09, 2.08401e-08, -3.273556e-09, -1.453651e-08, 8.356608e-09, 
    -2.858961e-09, 6.629399e-08, -4.573337e-09, 2.403706e-08, -3.241104e-08, 
    -1.691416e-08, -1.337327e-08, 7.632542e-08, 5.071286e-09, -2.188295e-08, 
    -3.344582e-08, 2.232667e-08, 3.055032e-08, -6.59507e-08, 2.887731e-08, 
    -5.698831e-08, 5.192504e-08, -7.670775e-08, 5.039391e-08, 3.239728e-08, 
    -1.019913e-08, 6.608369e-08, 6.914433e-10, -3.703332e-08, -8.747769e-08, 
    1.65309e-07, 4.256771e-08, -9.00132e-08, 2.208225e-08, 7.270199e-08, 
    -2.759685e-08, -5.877024e-08, -5.548861e-08, -3.792877e-09, 7.051156e-09, 
    3.160326e-08, -6.823171e-08, 9.920393e-09, 1.879315e-08, -2.183689e-08, 
    -2.230479e-09, -8.013063e-08, 1.094115e-07, -2.477086e-07, -4.092101e-09, 
    -3.799983e-10, 4.384623e-08, 1.66778e-08, 2.372188e-08, 5.634319e-08, 
    5.065584e-08, 1.498341e-08, 1.907091e-08, -1.971426e-08, 5.774325e-09, 
    -1.561426e-08, -1.21951e-07, -4.499299e-08, 2.811191e-09, -2.399381e-08, 
    4.788888e-09, 3.046836e-09, 4.692879e-09, -1.55839e-08, -4.986629e-08, 
    -3.894951e-08, 2.498826e-08, -1.121346e-07, 6.942236e-08, 3.148159e-09, 
    4.899846e-09, 7.308762e-08, 3.080174e-09, -4.483833e-08, -8.307268e-09, 
    1.368852e-08, -1.578577e-09, -6.104813e-09, 4.941138e-08, -1.049321e-07, 
    3.124919e-07, -1.7068e-08, -8.316022e-09, -6.290503e-08, 9.586245e-09, 
    1.067741e-08, 9.193272e-09, 8.687095e-10, -5.84896e-09, 5.626083e-08, 
    3.053646e-08, 1.472653e-07, 2.398878e-08, -1.05893e-08, -4.919076e-08, 
    -9.554526e-09, -9.50655e-09, -2.138734e-09, 5.141771e-09, 1.971728e-09, 
    3.701768e-09, 5.788905e-09, -1.487891e-09, 6.416911e-10, 5.332384e-08,
  -5.031802e-08, -5.643142e-08, 2.038996e-08, -7.208496e-08, 2.146203e-08, 
    -1.020271e-08, 3.774403e-09, 4.272124e-09, 7.15977e-09, 1.427884e-08, 
    -2.127763e-09, -4.905451e-08, -5.061338e-10, -1.584385e-08, 1.289322e-08, 
    -1.32206e-08, 6.057674e-08, -4.475282e-09, 2.434425e-08, -2.494357e-08, 
    -1.8538e-08, -1.256535e-08, 7.769904e-08, 5.375568e-09, -2.175534e-08, 
    -3.784021e-08, 7.868152e-08, 2.216007e-08, -2.496336e-09, 8.757297e-09, 
    -8.304096e-08, 5.794709e-08, -4.146023e-08, 1.004837e-07, 3.245759e-08, 
    -3.340301e-08, 5.629895e-08, 8.564314e-10, -6.32665e-08, -8.807329e-08, 
    1.610485e-07, 4.396088e-08, -9.896274e-08, 1.773399e-08, 5.03926e-08, 
    3.868308e-09, -5.852473e-08, -5.507735e-08, 1.123408e-08, 7.48679e-09, 
    3.08826e-08, -7.001131e-08, 9.534392e-09, 1.876229e-08, -2.175321e-08, 
    4.712888e-09, -8.672714e-08, 1.166933e-07, -2.781144e-07, -3.639713e-09, 
    -4.025651e-09, 4.363642e-08, 1.757644e-08, 3.257223e-08, 4.798717e-08, 
    4.876347e-08, 2.343199e-08, 2.180195e-08, 3.260993e-09, -1.299668e-09, 
    -1.526428e-08, -1.115259e-07, -4.405069e-08, 3.816922e-09, -2.444199e-08, 
    5.729817e-09, 4.146472e-09, 5.986692e-09, -2.091537e-08, -4.997196e-08, 
    -3.60194e-08, 2.774692e-08, -1.145556e-07, 7.342715e-08, 3.178002e-09, 
    5.519496e-09, 5.727702e-08, 2.610932e-09, -4.251018e-08, -1.159469e-08, 
    1.463991e-08, -1.419311e-09, -6.606058e-09, 4.957553e-08, -1.263259e-07, 
    3.109041e-07, -1.612861e-08, 4.533103e-08, -6.379105e-08, 1.031194e-08, 
    2.73053e-08, 7.269421e-09, -2.580862e-09, -5.554952e-09, 7.86647e-08, 
    2.978391e-08, 3.166426e-07, 5.321886e-08, 2.11694e-08, -3.580294e-08, 
    -2.837169e-09, -6.422852e-09, -1.223952e-09, 5.595666e-09, 3.214154e-09, 
    3.943117e-10, 2.2508e-09, -6.638203e-09, 1.033271e-10, 5.744801e-08,
  -4.47983e-08, -5.663446e-08, 1.341073e-08, -7.711947e-08, 2.200159e-08, 
    2.534762e-09, 2.600245e-09, 1.239914e-08, 6.886921e-09, 2.086449e-08, 
    -2.854222e-09, -6.307368e-08, 4.135245e-09, -1.581816e-08, 1.560556e-08, 
    -1.514557e-08, 5.745433e-08, -4.192543e-09, 2.531931e-08, -1.563967e-08, 
    -1.970898e-08, -1.213834e-08, 7.894869e-08, 5.698666e-09, -2.145111e-08, 
    -4.088724e-08, 6.823143e-08, 1.034186e-08, -1.664557e-08, 3.768992e-08, 
    -6.952064e-08, 5.683228e-08, -2.910701e-08, 8.909046e-08, 3.26238e-08, 
    -4.65609e-08, 4.534886e-08, 3.342109e-10, -6.969435e-08, -8.484196e-08, 
    1.647979e-07, 4.330059e-08, -1.037085e-07, 1.726134e-08, 5.698416e-08, 
    2.619322e-08, -5.870936e-08, -5.402853e-08, 1.970739e-08, 8.211146e-09, 
    2.985084e-08, -7.157996e-08, 1.126559e-08, 1.839999e-08, -2.17426e-08, 
    -3.044079e-09, -8.926395e-08, 1.206503e-07, -2.982281e-07, -2.476185e-09, 
    -5.924448e-09, 4.345111e-08, 1.833541e-08, 3.238406e-08, 3.759182e-08, 
    5.060838e-08, -3.085074e-08, 3.125433e-08, 4.871117e-08, -6.35805e-09, 
    -1.519743e-08, -9.911514e-08, -4.518211e-08, 4.57112e-09, -2.51189e-08, 
    2.605248e-09, 4.190753e-09, 6.08668e-09, -1.696741e-08, -5.015249e-08, 
    -5.584218e-08, 2.964697e-08, -1.160173e-07, 7.550011e-08, 4.285539e-09, 
    5.249149e-09, 5.280663e-08, 2.428806e-09, -4.032385e-08, -1.423268e-08, 
    1.515514e-08, -3.385958e-09, -6.862479e-09, 4.837868e-08, -1.339083e-07, 
    3.089134e-07, -1.495819e-08, 7.756034e-08, -6.556957e-08, 1.277654e-08, 
    3.4918e-08, 7.556977e-09, 2.107356e-09, -5.365109e-09, 6.529012e-08, 
    2.9484e-08, 3.117616e-07, 7.062681e-08, 4.478943e-08, -2.657384e-08, 
    3.980404e-09, -2.320576e-09, 2.137313e-10, 5.756192e-09, 3.741661e-09, 
    1.118201e-09, -8.586198e-11, 7.281002e-10, 3.368115e-10, 6.196547e-08,
  -4.285835e-08, -5.302763e-08, 9.111545e-09, -8.026814e-08, 2.032039e-08, 
    1.073954e-08, 1.737135e-09, 1.407898e-08, 7.592462e-09, 2.083721e-08, 
    -2.66823e-09, -7.233257e-08, 4.482217e-09, -1.597959e-08, 1.521857e-08, 
    1.265903e-10, 5.636221e-08, -4.312142e-09, 2.454138e-08, -1.05008e-08, 
    -2.016009e-08, -1.226067e-08, 7.996277e-08, 6.262098e-09, -1.996818e-08, 
    -4.16419e-08, 6.282471e-08, -8.854386e-09, -2.778438e-08, 3.156356e-08, 
    -7.596941e-08, 4.032063e-08, -1.250623e-08, 1.113231e-07, 3.248647e-08, 
    -6.181335e-08, 3.611726e-08, -1.08605e-09, -7.40722e-08, -8.23246e-08, 
    1.781403e-07, 4.108188e-08, -1.052003e-07, 4.241169e-09, 5.740162e-08, 
    3.883292e-08, -5.967445e-08, -5.22935e-08, 2.782262e-08, 1.103706e-08, 
    2.922027e-08, -7.288736e-08, 1.455608e-08, 1.886633e-08, -2.184532e-08, 
    -3.290893e-09, -9.110181e-08, 1.215745e-07, -3.124838e-07, -1.178677e-09, 
    -5.740276e-09, 4.303683e-08, 1.873491e-08, 3.430718e-08, 2.731135e-08, 
    2.700062e-08, -3.50658e-08, 7.906465e-09, 3.76408e-08, -6.734581e-09, 
    -1.556873e-08, -1.299802e-07, -4.142066e-08, 5.158199e-09, -2.55196e-08, 
    -1.910098e-08, 3.74834e-09, 5.671609e-09, -1.22781e-08, -4.944422e-08, 
    -6.082951e-08, 3.003861e-08, -1.168613e-07, 7.58962e-08, 4.365347e-09, 
    4.116373e-09, 5.087441e-08, 2.203706e-09, -3.847997e-08, -1.634282e-08, 
    1.494891e-08, -2.908019e-09, -7.056656e-09, 4.618967e-08, -1.502733e-07, 
    3.003138e-07, -1.50666e-08, 8.855091e-08, -6.697655e-08, 1.419757e-08, 
    3.974992e-08, 7.522345e-09, 5.231215e-09, -6.860219e-09, 5.710285e-08, 
    2.93212e-08, -2.626894e-08, 8.062102e-08, 6.160212e-08, -2.100683e-08, 
    1.156968e-08, -1.437229e-09, 2.835577e-09, 6.568371e-09, 3.40151e-09, 
    3.728064e-09, 8.244768e-09, -8.465406e-10, 7.114949e-10, 6.575237e-08,
  -4.066828e-08, -5.452148e-08, 4.353979e-09, -8.030247e-08, 1.770218e-08, 
    1.325566e-08, 9.652013e-10, 1.335889e-08, 6.946266e-09, 1.907301e-08, 
    -2.599791e-09, -7.683229e-08, 4.808498e-09, -1.617263e-08, 1.449325e-08, 
    6.150088e-09, 5.756402e-08, -4.203116e-09, 2.350791e-08, -6.34418e-09, 
    -2.091224e-08, -1.288936e-08, 8.04655e-08, 7.314384e-09, -1.744729e-08, 
    -3.956188e-08, 6.121059e-08, -1.872831e-08, -3.039008e-08, 4.099957e-08, 
    -7.974336e-08, 7.886251e-08, -5.3044e-09, 1.054052e-07, 3.213609e-08, 
    -7.434483e-08, 3.05789e-08, -1.069651e-09, -7.784388e-08, -8.044067e-08, 
    1.723484e-07, 3.910145e-08, -1.103292e-07, 2.730374e-09, 5.399011e-08, 
    6.386131e-08, -6.060827e-08, -5.106892e-08, 3.50456e-08, 9.447319e-09, 
    2.881427e-08, -7.411245e-08, 1.87106e-08, 2.12181e-08, -2.198058e-08, 
    -7.185008e-11, -9.200699e-08, 1.19339e-07, -3.186122e-07, -4.251604e-10, 
    -5.515858e-09, 4.306912e-08, 1.886997e-08, 3.580089e-08, 1.961889e-08, 
    5.246648e-09, -4.008825e-08, 7.689778e-10, 4.346271e-08, -6.468554e-09, 
    -1.595549e-08, -1.669555e-07, -4.008393e-08, 5.580205e-09, -2.574275e-08, 
    -8.198413e-09, 4.119954e-09, 5.924392e-09, -1.129272e-08, -4.778667e-08, 
    -6.090238e-08, 2.9852e-08, -1.216076e-07, 7.486915e-08, 2.272827e-09, 
    1.911985e-09, 4.918707e-08, 1.854005e-09, -3.694437e-08, -1.806939e-08, 
    1.534613e-08, -1.863828e-09, -7.341157e-09, 4.273031e-08, -1.658639e-07, 
    2.806125e-07, -1.961403e-08, 9.401333e-08, -6.77901e-08, 1.564904e-08, 
    4.253161e-08, 7.643592e-09, 7.580311e-09, -7.014123e-09, 5.228685e-08, 
    2.938486e-08, -1.689955e-08, 8.845996e-08, 7.974791e-08, -1.719786e-08, 
    1.848321e-08, -2.846946e-09, 7.136805e-09, 1.822423e-08, 2.681418e-09, 
    9.132009e-10, 3.541743e-09, -4.100968e-09, 5.179004e-10, 6.513937e-08,
  -3.899083e-08, -5.327763e-08, -3.46779e-09, -8.272411e-08, 1.366755e-08, 
    1.214005e-08, -5.965148e-10, 1.05191e-08, 4.212438e-09, 1.606202e-08, 
    -2.996217e-09, -7.788083e-08, 3.022819e-09, -1.635374e-08, 1.394767e-08, 
    -1.766131e-08, 9.137288e-08, -5.432526e-09, 2.073696e-08, -5.297238e-09, 
    -2.281706e-08, -1.402498e-08, 7.974825e-08, 9.705559e-09, -1.252204e-08, 
    -3.780758e-08, 3.88244e-08, -2.44969e-08, -3.844218e-08, 5.154868e-08, 
    -8.285735e-08, 7.970868e-08, -2.664024e-09, 7.83383e-08, 3.117941e-08, 
    -8.778773e-08, 2.783838e-08, -5.022969e-10, -8.104973e-08, -7.944871e-08, 
    1.663358e-07, 3.603134e-08, -1.034302e-07, 1.807972e-09, 6.002472e-08, 
    6.595599e-08, -6.052358e-08, -4.919957e-08, 4.103947e-08, 5.173007e-09, 
    2.714501e-08, -7.57683e-08, 2.464976e-08, 1.924098e-08, -2.229072e-08, 
    2.632873e-09, -9.324356e-08, 1.106275e-07, -3.116048e-07, -7.250378e-11, 
    -5.170818e-09, 4.112792e-08, 1.925616e-08, 3.75316e-08, 2.899831e-08, 
    -2.742695e-09, -4.283959e-08, 7.47491e-10, 4.202172e-08, -6.840423e-09, 
    -1.655155e-08, -1.769432e-07, -3.350544e-08, 6.452069e-09, -2.442673e-08, 
    -9.017981e-09, 3.529891e-09, 5.364484e-09, 1.255452e-08, -4.427932e-08, 
    -5.806828e-08, 2.833529e-08, -1.184181e-07, 7.058463e-08, 1.217586e-10, 
    -2.646289e-09, 4.708238e-08, 1.115609e-09, -3.510033e-08, -1.958995e-08, 
    1.553337e-08, -1.429886e-09, -7.662891e-09, 3.915133e-08, -1.866441e-07, 
    2.581489e-07, -2.359109e-08, 9.158032e-08, -6.693006e-08, 1.468459e-08, 
    4.533797e-08, 7.85775e-09, 6.734183e-09, -6.542336e-09, 5.034883e-08, 
    2.990225e-08, -1.810884e-08, 1.130592e-07, 1.043103e-07, -9.789005e-09, 
    2.66599e-08, -3.601258e-09, 8.355983e-11, 5.529159e-09, 1.595367e-09, 
    1.23714e-09, -5.827573e-08, 4.693845e-10, 1.186467e-08, 5.88044e-08,
  1.014325e-13, 2.511474e-13, 1.757199e-13, 1.932445e-13, 3.385492e-13, 
    5.449525e-13, 2.906692e-13, -1.344813e-14, -3.004398e-13, -4.223394e-13, 
    2.596515e-13, 4.371814e-13, -1.954593e-13, -1.363365e-13, 1.114148e-14, 
    2.051239e-13, 3.868557e-13, -2.406585e-12, 3.928098e-13, -2.996165e-13, 
    -9.564255e-13, -1.959203e-12, -5.899413e-13, 6.506361e-13, -1.253807e-12, 
    -4.897595e-13, -1.464946e-13, 2.331721e-13, 3.025305e-14, -5.640697e-15, 
    8.441095e-14, -7.094287e-15, -6.57393e-14, -2.213618e-14, -5.084854e-14, 
    1.048529e-13, -7.20533e-13, -3.081145e-12, 1.641134e-13, 2.002351e-12, 
    -1.938353e-13, 5.36458e-14, 2.699935e-13, 2.553144e-13, 1.728682e-13, 
    1.440271e-13, 3.268521e-13, 2.949692e-12, 8.06412e-13, 9.685632e-12, 
    -9.272626e-13, -4.30602e-13, 1.799453e-12, 1.471284e-12, 1.79115e-13, 
    -1.308932e-12, 1.016597e-13, 1.911241e-12, 2.483538e-13, 1.993149e-13, 
    1.056471e-12, 1.111049e-13, 1.737741e-13, -1.774714e-12, -4.765347e-12, 
    -2.16225e-14, -8.665041e-14, 1.495908e-13, 1.103926e-13, 3.271102e-14, 
    1.431424e-13, 1.884638e-13, 1.050323e-13, -2.269837e-13, -1.05587e-13, 
    1.707925e-13, -1.199169e-14, -4.465801e-13, -1.93967e-12, -8.190753e-13, 
    -1.940956e-13, -1.927487e-12, 1.277929e-12, -1.085854e-12, 2.441318e-13, 
    3.539213e-13, 3.655734e-13, -8.280323e-16, 2.22206e-12, 1.4817e-12, 
    5.781723e-13, 5.382963e-13, -1.215822e-12, -6.492457e-13, 1.052024e-13, 
    3.336409e-13, 4.697357e-14, 5.584343e-13, 8.884162e-13, -2.55013e-14, 
    -4.090775e-12, -1.487137e-13, 1.090296e-12, -1.337785e-12, -3.53748e-13, 
    -2.203339e-13, -7.089462e-13, -1.081984e-12, -1.197324e-12, 
    -5.628818e-13, -3.376569e-13, -4.61156e-14, 8.539415e-14, 6.094031e-14, 
    7.778504e-13, 9.861924e-13, 6.526693e-13, -3.541503e-13, 1.060386e-13, 
    -3.762342e-13,
  5.394586e-13, 5.674487e-13, 4.96407e-13, 4.142744e-13, 3.468544e-13, 
    2.527921e-13, 2.625867e-13, 2.008408e-13, 1.172826e-13, 3.961799e-14, 
    1.389765e-13, -1.295718e-13, -2.909888e-13, -3.774737e-13, -4.403153e-13, 
    1.460057e-13, -1.309991e-13, -1.980719e-14, -3.121037e-13, -5.913065e-13, 
    -1.014586e-12, -2.242789e-12, -2.829391e-12, 1.721395e-13, 5.633631e-14, 
    -9.013974e-14, -2.290729e-13, -3.774787e-14, 6.237652e-16, -1.41719e-13, 
    7.854504e-14, 2.278273e-13, 8.989601e-14, 3.193112e-14, 1.436278e-13, 
    1.177311e-13, -7.5304e-13, 7.045264e-16, 4.309305e-13, 2.344901e-13, 
    -6.785499e-13, 3.749734e-13, -4.282836e-13, 3.972859e-13, -3.552281e-13, 
    -7.450214e-13, -5.260494e-13, 7.409535e-13, -5.966863e-13, 4.336238e-13, 
    8.150444e-14, -2.876453e-13, 8.370708e-13, 1.755985e-12, 6.218614e-13, 
    -1.027331e-12, 6.50396e-13, -1.374107e-12, -2.75925e-13, 2.284507e-13, 
    7.794117e-13, 1.613967e-13, 8.252883e-14, -2.558691e-13, -1.935991e-13, 
    1.085282e-13, -1.710885e-13, -9.017412e-14, -1.597188e-13, 6.035411e-15, 
    -1.87764e-12, 3.022736e-13, 5.973812e-13, 7.695199e-14, 3.027559e-12, 
    -1.441909e-13, -4.372342e-13, 5.599151e-13, -2.101229e-12, 3.835319e-13, 
    2.054183e-13, 1.26563e-12, -1.471267e-12, 3.289569e-13, 5.438472e-13, 
    9.874534e-13, -7.858476e-13, 2.012404e-13, 2.804411e-13, 1.317616e-13, 
    3.584255e-13, 1.864344e-14, -1.384029e-14, -3.901852e-14, 1.547339e-13, 
    1.511654e-13, 2.010112e-13, -1.508592e-13, 3.148185e-13, -2.59716e-13, 
    2.571746e-13, -4.717423e-13, -1.703766e-12, -8.017756e-13, -1.641695e-14, 
    1.200354e-13, -4.679596e-14, -3.3139e-13, -7.914433e-13, -6.059612e-13, 
    -6.824912e-13, -1.967533e-13, 6.1938e-14, 1.482574e-13, -4.535736e-14, 
    1.130546e-12, -3.985687e-13, -1.489988e-12, -3.543925e-13, -6.269579e-15,
  1.901118e-13, 1.687539e-14, -7.92838e-14, -1.434963e-14, 1.17642e-13, 
    2.048778e-13, 3.54286e-13, 1.682682e-13, 1.035422e-13, -1.494915e-13, 
    -3.934353e-14, -6.827872e-15, 3.450018e-14, 3.538836e-15, -7.009671e-14, 
    1.413175e-13, 1.508099e-13, -4.394402e-14, 3.386787e-13, 4.688333e-13, 
    5.441064e-13, 3.900907e-13, 5.225959e-13, 2.378653e-13, 7.649437e-13, 
    8.316126e-13, 6.576545e-13, 3.436834e-13, 2.090411e-13, 1.905698e-13, 
    2.326611e-13, 2.137179e-15, 1.077471e-13, 7.373269e-14, 7.042977e-14, 
    1.751377e-13, -1.808149e-12, 3.041664e-14, -3.312906e-13, 1.621341e-12, 
    -2.230161e-13, -1.055545e-12, 4.277759e-13, 1.626431e-13, -2.222528e-13, 
    -1.428163e-13, -8.001377e-13, 7.332746e-13, -4.173967e-13, -3.679513e-13, 
    5.25394e-13, -6.284695e-13, 1.602192e-12, -2.11523e-11, 1.17962e-17, 
    -1.737679e-12, -5.998813e-13, -9.505785e-13, 9.290873e-13, -5.518364e-13, 
    1.378522e-12, -3.040068e-13, -2.081529e-13, -1.089406e-14, -2.421896e-13, 
    -2.216699e-13, 1.185579e-13, -2.804701e-14, -3.441691e-15, 2.297051e-13, 
    -6.360606e-13, 1.095096e-13, 1.036685e-12, 3.943235e-13, -1.365782e-13, 
    -3.188241e-12, -9.286669e-14, 5.815314e-13, -3.711944e-12, -1.099953e-13, 
    1.797389e-12, 1.198585e-12, -3.065881e-13, 3.097661e-13, 6.867701e-13, 
    3.707173e-13, 1.675285e-12, 5.116463e-13, 3.578787e-13, 1.449278e-12, 
    -4.421463e-14, -2.131545e-13, 3.659018e-13, -8.130718e-13, -3.051726e-14, 
    -2.675388e-13, 3.871348e-13, -1.391942e-13, 6.982193e-13, 1.32705e-12, 
    -4.402312e-13, 2.668447e-13, 2.830947e-13, 8.176619e-14, -3.093081e-13, 
    -8.126694e-13, -7.995271e-13, -1.183303e-12, -2.10533e-12, -2.294234e-12, 
    -7.767675e-13, -4.718448e-14, 1.706968e-13, 4.386769e-13, 1.228323e-13, 
    3.56673e-13, 1.709329e-12, 1.296913e-11, -5.398086e-13, -4.498485e-13,
  2.768341e-13, 2.345901e-13, 2.674527e-13, 3.551465e-13, 4.295592e-13, 
    4.504591e-13, 3.288064e-13, 5.67324e-14, -2.902262e-13, -5.628692e-13, 
    -3.878287e-13, -3.282097e-13, -5.56083e-13, -4.018591e-13, -6.833423e-13, 
    -1.06247e-13, 2.135639e-13, -1.87593e-13, -1.39961e-13, 2.476491e-13, 
    8.844314e-14, -1.235401e-13, -2.722544e-13, -5.982437e-13, -2.171374e-12, 
    -2.649811e-12, -1.526557e-16, 2.211981e-13, 6.362966e-14, 4.977962e-13, 
    1.623701e-14, -2.640943e-13, -7.940593e-13, 7.921441e-14, 8.01581e-14, 
    1.985495e-13, -1.027194e-12, 3.617662e-13, 2.009504e-13, -1.057945e-13, 
    -1.559308e-14, 2.806505e-13, 3.041942e-13, 4.110839e-14, 1.506711e-13, 
    -7.177731e-13, -7.858228e-13, 3.803555e-13, 1.340245e-12, 6.992019e-12, 
    -5.490088e-13, -2.505912e-13, 6.456336e-13, 2.360034e-12, 1.304571e-13, 
    -1.432632e-12, 2.071218e-12, -1.16586e-12, -1.28289e-13, -1.51938e-12, 
    3.367168e-13, 5.426076e-13, -1.85936e-12, 3.503753e-13, -7.660262e-14, 
    -1.169481e-13, -2.668699e-14, -4.135026e-13, -2.355338e-13, 3.195916e-13, 
    1.177392e-13, 4.973799e-14, -2.405021e-14, 4.711231e-13, -4.889048e-13, 
    -2.535944e-12, 2.112739e-12, 2.124172e-12, -2.414654e-11, -1.790651e-13, 
    1.183595e-12, 4.944895e-13, -2.548378e-13, -1.947956e-12, -2.516876e-13, 
    1.654371e-13, -9.672818e-15, -4.719697e-13, -2.726049e-13, -3.26697e-13, 
    -3.011064e-13, -3.71728e-12, 4.544559e-13, -1.224042e-12, -5.813405e-13, 
    -1.433933e-12, -5.940636e-13, -5.928591e-14, -4.792847e-12, 
    -2.138728e-12, 4.824474e-13, -1.849837e-12, 3.692532e-13, 3.719984e-13, 
    -3.288619e-13, -2.648159e-13, -6.122186e-13, -2.619016e-13, 
    -3.702594e-14, 9.0844e-14, 2.871869e-13, 2.049055e-13, 2.103179e-13, 
    2.589595e-13, 1.437461e-13, 5.523804e-13, 5.523066e-12, 3.765992e-12, 
    -2.139781e-15, -6.733225e-13,
  7.978895e-13, 5.653811e-13, 4.660439e-13, 3.891054e-13, 4.021228e-13, 
    5.602463e-13, 8.123502e-13, 4.889977e-13, -7.424616e-14, -8.920364e-13, 
    -6.107614e-13, -4.475864e-13, -9.300893e-14, 2.224054e-13, 3.629319e-13, 
    -1.628503e-13, 3.219647e-14, -9.222206e-13, -3.109978e-13, 1.351419e-13, 
    6.94278e-13, 1.515177e-13, -8.126e-13, -1.549538e-12, -2.028183e-12, 
    -2.39983e-12, 1.192435e-12, 2.987333e-13, -3.241851e-14, -3.89716e-13, 
    4.360401e-13, 4.325984e-13, 6.79734e-13, -6.76903e-13, -9.925949e-13, 
    -2.866873e-13, -1.015052e-12, 1.282651e-12, 1.840195e-13, 9.427847e-13, 
    2.261413e-13, 3.993472e-13, 8.790191e-14, 2.28258e-13, -2.204847e-12, 
    -1.224326e-12, -1.076916e-13, -1.405001e-12, 3.231243e-12, 2.729719e-11, 
    -3.912703e-13, -6.483425e-13, -9.578449e-13, -1.205763e-12, 8.855832e-14, 
    -1.427428e-12, 5.736051e-12, -5.887485e-13, 5.22915e-14, -1.566768e-12, 
    -2.989831e-13, -1.739997e-13, -3.622103e-14, 9.406365e-14, 1.724565e-13, 
    1.835476e-13, -7.121803e-13, -2.41307e-13, 4.791167e-13, -1.831785e-12, 
    1.416645e-13, -5.916378e-13, -1.980083e-13, 4.49446e-13, -1.311479e-13, 
    -1.214806e-12, 7.576231e-13, -7.206596e-13, -4.679602e-12, 1.023431e-12, 
    2.05766e-13, 5.907754e-13, -7.820133e-13, -2.359418e-12, -1.874167e-12, 
    -2.745582e-13, -3.095579e-13, -5.700995e-14, 1.266357e-13, -4.014844e-14, 
    -4.889422e-13, 2.430722e-13, 6.50105e-14, 1.687017e-12, 5.364043e-13, 
    8.373915e-12, -4.791334e-13, -3.971823e-13, -3.650635e-12, 4.32332e-13, 
    3.114176e-13, 1.075504e-12, 6.272257e-13, 1.396364e-12, -5.176415e-14, 
    -2.349787e-13, -2.632616e-13, 5.531686e-14, 3.041734e-13, 2.793321e-13, 
    7.308321e-13, 9.107992e-13, 3.050338e-14, 9.361956e-14, -9.242607e-15, 
    1.969541e-12, 7.251203e-12, -1.64157e-11, -1.00828e-12, 5.892509e-14,
  4.303502e-14, 6.257495e-14, -3.720635e-14, 8.056056e-14, 5.290074e-13, 
    6.546153e-14, -8.285039e-15, 2.583073e-13, 3.062689e-13, 9.316853e-13, 
    -2.807476e-14, 3.285566e-13, -6.281781e-13, -1.747255e-12, -9.202777e-13, 
    -7.097656e-14, -4.333617e-13, 1.999928e-13, -6.445885e-13, -6.743356e-13, 
    -9.787865e-13, 1.631043e-12, 1.673897e-12, 3.159834e-13, -1.71603e-12, 
    -1.256481e-12, -5.119377e-13, -1.658534e-13, 7.643469e-13, -9.849205e-13, 
    -3.03034e-12, -1.759856e-12, -1.945569e-12, 1.593711e-12, -2.413583e-12, 
    3.506501e-13, -6.867479e-13, 6.141719e-13, 1.058612e-12, -7.319173e-13, 
    1.690284e-12, -8.886364e-13, 1.28321e-13, -2.345997e-14, 7.907147e-13, 
    -2.93289e-12, -4.359152e-13, 3.36408e-12, 2.629344e-12, 1.508383e-11, 
    -8.927824e-13, -5.036124e-12, 4.221682e-12, 2.794617e-12, 3.18176e-13, 
    -1.313685e-12, -4.037701e-12, -1.096262e-13, 1.136882e-12, -4.458343e-13, 
    1.091141e-12, -2.026726e-12, 6.035311e-13, -1.512651e-13, 2.742168e-13, 
    -3.485684e-13, 2.486802e-12, -1.287345e-12, 2.421771e-12, -4.379136e-13, 
    -2.527936e-12, -1.853143e-12, 7.23463e-13, -1.207714e-12, -4.977785e-12, 
    -1.901548e-12, -2.697911e-13, -8.499451e-14, -6.340979e-12, 3.000669e-12, 
    1.551648e-12, -3.703225e-13, -1.206757e-12, -1.379133e-12, -1.245629e-12, 
    -4.563003e-12, -3.512954e-12, -4.79769e-13, 6.242398e-13, -2.436218e-12, 
    -7.524953e-13, -3.021666e-13, 3.215345e-13, 3.01334e-12, 2.382955e-13, 
    -2.644374e-12, 5.095119e-13, -5.669493e-13, 4.331105e-12, 2.699979e-13, 
    -2.306391e-12, 7.383018e-13, 5.563692e-13, -1.716792e-12, -3.943373e-13, 
    -8.583551e-13, -1.037295e-12, 1.302694e-12, 1.467063e-12, 8.031215e-13, 
    5.489637e-13, 1.102521e-12, 1.269401e-13, 2.167475e-12, -7.22436e-13, 
    1.702241e-12, 2.549211e-12, -2.406003e-12, -2.191997e-13, 9.322126e-13,
  -8.20996e-13, -1.009609e-13, 7.822909e-14, -4.905798e-14, 1.357539e-12, 
    4.307249e-13, 5.371398e-13, 2.517e-12, 4.099124e-12, -4.486564e-12, 
    -4.715048e-12, -2.075548e-12, -6.054365e-12, -5.841647e-12, 
    -3.173004e-12, -7.503748e-13, -9.559492e-13, 1.170161e-12, -4.239109e-13, 
    -1.494291e-12, -8.770623e-13, 7.766704e-13, 2.02173e-12, 2.031056e-12, 
    1.888767e-14, 6.67684e-12, 2.360348e-12, -8.492582e-12, 2.303172e-12, 
    2.830639e-12, 1.632722e-13, 3.580428e-12, -3.281306e-12, 3.723272e-13, 
    -1.371389e-12, 3.624614e-12, -4.575812e-13, 6.891085e-13, 2.985528e-13, 
    -1.856765e-13, -5.719286e-13, 6.60956e-12, -1.154979e-12, 5.790255e-13, 
    -6.486797e-12, 2.668712e-12, 2.490647e-13, 2.061129e-13, -1.505537e-12, 
    -9.481041e-12, 2.47713e-12, -4.142339e-12, 1.308592e-13, 1.280222e-11, 
    2.166059e-13, -8.486961e-13, -7.86135e-13, -4.300033e-13, 1.676712e-12, 
    -9.793971e-13, 3.728198e-12, 7.861767e-14, -5.039677e-12, -1.226527e-12, 
    -1.382866e-13, 1.890101e-11, 1.576513e-11, -3.721731e-12, -8.734e-12, 
    2.989234e-12, -5.286424e-12, -1.139186e-12, -2.305919e-12, -6.473572e-13, 
    -3.291759e-12, -1.542252e-12, -3.152756e-13, -1.955519e-13, -1.75935e-11, 
    2.345804e-12, 3.511788e-12, 3.118614e-12, -7.677609e-13, 7.080184e-12, 
    2.369174e-12, -4.857212e-12, -3.569631e-12, 6.522144e-13, -1.419718e-12, 
    1.842235e-12, -1.883813e-12, -1.562059e-12, -2.083195e-13, 7.355977e-13, 
    3.070169e-12, -7.35825e-12, -1.112485e-12, -8.293227e-13, 1.361029e-11, 
    2.755832e-12, -6.517425e-13, 1.196876e-12, 7.458097e-13, -9.829897e-12, 
    -1.583164e-12, 4.419382e-13, -1.595807e-13, 1.916592e-12, 1.467507e-12, 
    9.766771e-13, 1.078929e-12, 2.761472e-12, 3.55245e-12, 5.104944e-13, 
    1.062497e-12, -4.280937e-13, 9.904369e-13, -3.245246e-12, -1.213855e-13, 
    6.363146e-12,
  -1.511957e-12, 3.742173e-12, 6.394163e-12, 9.225565e-12, 1.267703e-11, 
    1.184081e-11, 1.373351e-11, 5.572376e-12, -8.245349e-12, 8.235634e-13, 
    -5.990985e-12, -1.486294e-11, -4.763412e-12, -1.57831e-11, -1.274464e-11, 
    2.119566e-12, 1.428124e-12, -5.984713e-12, 3.010717e-13, 3.628764e-13, 
    8.595347e-13, 1.06809e-12, 3.524958e-13, -7.326917e-13, 4.136136e-12, 
    1.779149e-11, 2.652406e-11, 4.849454e-13, 4.00957e-13, 9.286238e-12, 
    2.493616e-12, -5.900169e-12, -4.291678e-12, -6.515621e-12, 4.498568e-12, 
    1.859957e-12, -3.988404e-12, 5.130826e-13, 4.416689e-12, 3.699602e-12, 
    4.90511e-12, 3.736289e-12, 3.229222e-13, -4.289537e-14, -8.27366e-12, 
    1.18025e-11, 1.627559e-12, -3.201467e-13, 3.324119e-12, -2.505031e-11, 
    3.802937e-12, -3.701373e-12, 1.291234e-12, 5.253242e-12, -2.433942e-13, 
    -6.042944e-13, 5.943801e-12, 2.117084e-13, 1.53137e-12, 6.253498e-12, 
    -4.597434e-12, 9.369339e-12, -4.370837e-12, 2.440692e-12, -3.89544e-13, 
    1.087713e-11, -2.093159e-12, -2.624678e-12, -9.418633e-12, 9.775625e-12, 
    -2.902678e-12, 1.254769e-11, -7.827627e-13, -1.001477e-12, -5.923751e-12, 
    -5.633827e-13, -2.288308e-13, 3.516215e-13, -1.989688e-11, 3.350487e-12, 
    7.661038e-12, -3.124532e-11, 1.72623e-12, 2.276412e-11, 5.241918e-13, 
    -1.732836e-12, -2.011669e-12, 1.252665e-12, 6.988394e-13, 1.049466e-12, 
    8.915091e-14, -8.550271e-13, -4.315159e-13, 1.650557e-12, 8.426759e-12, 
    -1.834388e-12, 4.709177e-12, -5.011103e-12, 2.989775e-12, 7.295498e-13, 
    7.927714e-12, 2.561642e-12, 5.58234e-15, -4.279392e-11, -8.432699e-13, 
    1.372735e-12, -2.303713e-14, 1.365519e-12, 9.58178e-13, 2.127687e-12, 
    5.902889e-12, 3.584688e-12, -2.102263e-12, -8.054835e-12, -9.231504e-14, 
    -8.031964e-13, 1.667964e-12, -6.086437e-12, -2.999684e-14, 1.616574e-11,
  -4.60687e-12, 1.001421e-11, 1.186318e-11, 1.128136e-11, 1.123579e-11, 
    9.148293e-12, -9.512113e-12, 5.709655e-11, 4.864148e-11, 1.357908e-11, 
    1.092682e-12, -3.95517e-13, -2.345346e-13, -2.614853e-12, -1.495776e-11, 
    2.94782e-12, 3.006539e-13, -2.756823e-12, 1.075529e-13, 4.943268e-13, 
    6.777912e-14, -2.279288e-13, 7.727152e-14, -1.52986e-11, -6.712464e-12, 
    -1.558814e-11, 4.482748e-12, 2.828626e-12, -8.196999e-12, 1.468886e-11, 
    7.970569e-12, -1.231704e-11, 1.38739e-12, -4.876655e-12, -6.447509e-12, 
    1.184802e-11, -4.039957e-12, -5.114659e-14, 7.034262e-12, 2.584211e-13, 
    1.357459e-12, -4.452383e-12, -1.727229e-12, 2.004509e-12, 1.150968e-12, 
    8.798628e-12, 1.32222e-12, 7.017581e-13, 6.933276e-12, -1.036919e-11, 
    -2.452274e-13, -4.368728e-14, 4.818934e-12, -6.657008e-13, 1.850326e-14, 
    -7.158163e-14, 1.578737e-13, 5.153378e-13, -1.085132e-12, 1.840854e-11, 
    -2.501693e-11, 4.310885e-12, -5.372258e-12, -3.481337e-12, -6.35425e-12, 
    2.571277e-13, 9.532375e-13, 8.859025e-13, -5.742379e-11, 8.879175e-11, 
    1.463163e-12, -5.008022e-11, 5.714762e-12, -9.074907e-12, 5.002715e-12, 
    1.49436e-13, -3.868572e-13, 3.695239e-13, -4.272907e-12, 1.147116e-11, 
    9.673151e-12, -1.824281e-11, 1.15935e-12, -1.668504e-11, -1.025918e-11, 
    -4.777512e-12, 6.655954e-12, -2.31809e-12, 1.778301e-12, -3.278489e-13, 
    2.225664e-12, -1.473058e-11, -4.710399e-13, 2.259848e-12, 1.118494e-12, 
    -9.630074e-14, 7.015233e-12, -1.510003e-11, -3.143485e-12, 6.687539e-13, 
    -1.867173e-12, 2.305205e-13, -1.416749e-13, -4.227741e-11, 3.900213e-12, 
    4.810596e-13, -5.734302e-14, 1.488643e-12, 2.312317e-12, 1.128153e-12, 
    -2.754241e-12, -6.811773e-12, -4.648448e-12, 8.276491e-12, -7.082002e-12, 
    -5.801803e-13, 2.463307e-13, -3.942362e-12, -1.353223e-13, 5.350387e-12,
  -3.860468e-12, 3.595735e-12, 6.551926e-12, 7.931378e-12, 1.877054e-12, 
    2.250489e-11, 6.014911e-11, 3.898837e-11, -3.591238e-11, 1.617734e-11, 
    -8.437695e-15, 7.424839e-12, 9.954981e-12, 8.77437e-12, -2.209122e-12, 
    -1.378758e-12, -2.186401e-12, -4.336781e-12, -1.514205e-13, 4.826028e-12, 
    4.201861e-12, 1.217032e-11, 2.491723e-11, -1.635359e-11, -3.868572e-13, 
    -5.857259e-12, 1.066958e-11, 7.309037e-11, 1.155359e-11, -3.549022e-11, 
    7.526757e-12, 1.890238e-11, 8.965773e-12, 2.082834e-12, 7.850054e-12, 
    7.412848e-11, 2.518663e-12, -3.677961e-13, 3.615019e-11, -3.579587e-12, 
    2.140566e-12, 2.546297e-12, 5.595566e-12, 3.900991e-12, 1.221029e-11, 
    1.961875e-12, 1.29724e-12, 1.030731e-12, 5.316092e-12, 7.687288e-13, 
    -3.713557e-13, 7.310763e-12, 5.670048e-12, -4.054091e-13, -1.298679e-12, 
    5.83783e-13, 2.785217e-12, -2.895239e-13, -2.605444e-12, 2.044703e-11, 
    -3.896855e-11, 1.037226e-12, -9.41619e-12, -6.483569e-12, -7.063938e-12, 
    -5.81718e-12, 1.076572e-11, -8.338896e-11, -1.269601e-11, 1.576805e-11, 
    -3.570233e-11, 3.808243e-11, 2.328582e-11, 4.591827e-12, 2.770617e-12, 
    -3.179679e-13, -6.639828e-13, 5.767012e-12, 9.519104e-12, -1.151812e-11, 
    4.567818e-12, 4.750939e-11, -1.027789e-13, 1.877637e-11, -5.903611e-12, 
    5.28283e-12, 9.693468e-12, 5.034861e-14, 1.126559e-12, -1.421668e-12, 
    6.188716e-12, -8.724277e-12, -8.263945e-13, 1.119561e-11, -4.150125e-12, 
    -2.464462e-12, 1.979139e-12, 5.77669e-11, -8.635537e-12, -2.223444e-13, 
    -1.989653e-11, 1.050968e-12, -3.199489e-13, -2.246815e-11, -6.57141e-12, 
    1.434908e-12, 4.511391e-13, -4.162781e-12, 2.828071e-12, -2.004397e-12, 
    -1.131423e-11, -1.099948e-11, 1.697847e-11, 3.798523e-11, -1.138251e-11, 
    -4.987344e-13, 2.618045e-14, -3.029724e-12, 3.325028e-12, -7.49828e-12,
  1.54099e-12, 6.904921e-12, 1.253508e-11, 2.941558e-11, 9.048018e-11, 
    2.705025e-11, 1.495681e-11, -1.075835e-10, 5.812462e-12, -4.526024e-11, 
    1.352696e-12, -7.000178e-12, 5.983658e-12, 8.122725e-12, 7.042811e-12, 
    -3.414058e-12, -4.670719e-12, -7.159828e-12, 5.043535e-12, 7.419176e-12, 
    -8.325562e-13, -1.303202e-11, 1.895772e-11, -1.490275e-11, 2.407274e-11, 
    6.519008e-11, 2.592504e-11, -7.072898e-12, 4.952039e-12, -9.586998e-12, 
    1.750877e-11, 1.416045e-11, 8.291701e-12, -8.084755e-12, 4.164213e-11, 
    1.509015e-12, 1.018707e-12, -4.536649e-13, -5.151435e-13, -2.741296e-12, 
    1.649576e-11, 2.448763e-11, 2.278733e-12, 6.308738e-13, 2.488276e-11, 
    -2.214451e-11, 1.508571e-12, 1.004752e-13, -3.120371e-12, 7.278761e-13, 
    2.283618e-12, -2.049139e-11, 6.092959e-12, 1.63447e-13, 4.517026e-13, 
    3.805289e-13, 1.593803e-11, -1.276901e-12, -1.311673e-12, -1.737117e-11, 
    -2.473188e-11, -6.316059e-13, -1.454392e-14, -5.596523e-12, 
    -6.362399e-12, -1.081557e-11, 8.583245e-12, -1.22198e-10, 2.276035e-11, 
    1.373057e-11, -2.023459e-11, 2.938683e-11, 4.081713e-11, 3.988476e-12, 
    -1.188938e-13, -1.504463e-12, -7.601419e-13, -1.053843e-11, 3.317718e-12, 
    2.192468e-12, 6.579737e-13, 5.515033e-11, -8.276713e-14, 4.40048e-11, 
    -5.908385e-12, 7.188761e-11, 4.411527e-11, 7.387646e-12, 5.53519e-13, 
    -4.142298e-12, -1.35324e-11, -1.346634e-11, -9.730827e-13, -6.545875e-13, 
    -9.965917e-12, -4.869316e-12, -5.415957e-12, -1.262157e-11, 
    -1.883171e-11, -2.48821e-12, -2.70951e-11, -3.543832e-13, -7.156012e-13, 
    -2.328658e-12, -2.441236e-11, -1.260103e-13, 7.720491e-13, -9.778067e-12, 
    1.193523e-11, -4.511724e-12, -1.835332e-11, -7.639667e-12, 2.437328e-11, 
    2.764911e-11, -3.441358e-12, -1.164513e-13, 4.882206e-14, -2.071624e-12, 
    9.994165e-12, 2.715494e-12,
  -1.480738e-11, 2.832634e-11, 1.03797e-10, 8.121093e-11, 2.777989e-11, 
    -7.925438e-12, -2.448441e-11, 1.389417e-10, 1.641177e-10, 2.589295e-11, 
    -3.550582e-11, -2.193634e-11, -6.996737e-12, -2.146061e-13, 2.975198e-11, 
    -2.267675e-12, -5.111544e-12, -3.201384e-12, 5.244416e-14, -1.723288e-12, 
    5.828338e-12, -1.015477e-11, 4.531275e-11, -7.663314e-12, 4.736189e-11, 
    2.330338e-10, 2.41096e-12, -2.980005e-11, -5.199619e-12, 2.381972e-11, 
    4.613887e-11, 3.27377e-11, 6.49798e-11, -1.772027e-11, 6.217149e-11, 
    -8.992229e-11, -2.365108e-12, -3.606282e-13, 7.163803e-11, -2.278622e-13, 
    1.971772e-11, 2.931233e-11, -1.06426e-12, 1.197799e-12, 6.787937e-11, 
    1.699774e-11, 1.871003e-12, -4.378164e-13, -2.200085e-12, 3.996803e-15, 
    1.238844e-11, -7.264012e-11, 5.799516e-12, 1.082046e-12, 1.126257e-12, 
    -1.211253e-13, 1.569256e-11, -1.684253e-12, -3.27568e-12, -3.825078e-11, 
    -1.998945e-11, 3.047562e-13, 6.770695e-12, -4.077716e-12, -3.605494e-12, 
    -1.106142e-10, -1.017031e-11, -2.140169e-10, -1.441836e-11, 
    -4.063416e-14, -1.968981e-12, 6.057765e-11, -1.658925e-10, -9.796164e-12, 
    -1.059497e-12, -8.374412e-13, -5.729306e-13, -2.85256e-11, 1.568773e-13, 
    9.584444e-12, -4.707457e-12, 9.501486e-12, 6.930567e-13, 3.500999e-11, 
    -5.977585e-11, 2.464917e-12, 5.160072e-11, 2.189227e-11, -1.149875e-12, 
    -5.421441e-12, -6.476253e-11, -1.048337e-11, 2.692568e-13, -4.806553e-11, 
    -1.245559e-11, -3.482137e-12, -1.05379e-11, 9.922174e-12, -1.951239e-11, 
    -3.844702e-12, 3.894773e-12, -3.309575e-13, -2.002148e-13, 9.533416e-13, 
    4.254042e-12, -5.487832e-12, -1.798894e-11, 1.505063e-11, 1.014477e-11, 
    -7.849055e-12, -1.841938e-11, -6.012968e-12, 9.229284e-12, 1.381562e-11, 
    5.50715e-12, -8.988365e-14, 9.567347e-14, -1.357768e-13, 6.561925e-12, 
    -2.971523e-11,
  -4.297607e-11, 1.154794e-10, 1.142246e-10, 1.483746e-11, -3.271405e-11, 
    -6.088885e-11, -3.090483e-11, -2.12188e-11, 2.485079e-11, -2.086844e-10, 
    -4.632339e-11, 4.524114e-11, 7.060108e-11, -2.385625e-11, 4.312994e-11, 
    -1.089329e-12, -5.973067e-12, -3.462675e-12, -4.943379e-12, 9.384049e-12, 
    1.631206e-11, 5.701439e-12, 5.259437e-11, -3.568701e-12, 1.962031e-10, 
    4.375855e-10, -1.192246e-10, -2.207834e-11, -2.705725e-11, -7.12792e-11, 
    -2.855183e-11, 4.628586e-11, 1.669562e-10, -8.831602e-12, 9.47451e-11, 
    -2.613192e-10, -4.495071e-13, -2.537137e-13, 3.383491e-10, 1.161071e-13, 
    8.767475e-12, 3.040657e-11, 1.087597e-11, 9.700192e-13, 2.086331e-11, 
    3.559641e-11, 9.462431e-13, -1.759703e-13, 4.31184e-12, 1.491446e-13, 
    2.674858e-11, -9.006662e-11, 1.764988e-12, 2.618306e-12, 4.230116e-13, 
    -5.331291e-13, 3.839085e-11, -1.571987e-12, -8.80529e-12, -9.181406e-12, 
    -2.293654e-11, 2.15199e-11, -1.251887e-12, -3.5282e-12, -5.222667e-12, 
    -2.724345e-10, 3.086464e-11, -5.4785e-10, -5.717649e-13, 3.312661e-11, 
    -1.895506e-11, 9.461876e-11, -8.626055e-11, -3.785638e-11, -4.313283e-12, 
    -1.239009e-13, -2.109424e-13, -1.345396e-11, -1.248757e-12, 1.507061e-11, 
    -7.348122e-12, 7.815227e-12, 2.972067e-12, -9.490408e-12, -6.272161e-11, 
    -1.746965e-10, 1.466709e-10, 3.81617e-11, -1.78723e-12, -2.352785e-12, 
    -5.30942e-11, -1.33995e-12, 1.60516e-12, -5.189344e-11, -1.530398e-11, 
    -7.920354e-12, -1.518901e-11, 2.195177e-11, -4.638046e-11, -2.56497e-12, 
    1.613976e-11, 6.06562e-12, 3.538836e-14, 4.439643e-13, 6.783241e-12, 
    6.194156e-12, -4.207723e-11, -2.013878e-11, -8.200551e-12, -4.470202e-12, 
    -1.645972e-11, -5.430323e-12, -2.640999e-12, 2.077427e-11, 1.297851e-11, 
    -1.162848e-13, 1.48298e-13, 9.772738e-13, 2.293818e-12, -4.375789e-11,
  -2.557443e-11, 1.123148e-10, 1.104739e-11, -4.821321e-11, -4.729661e-11, 
    1.217915e-12, 1.784639e-11, -1.564209e-10, -2.375899e-11, -2.541125e-10, 
    5.589595e-11, -4.465317e-13, 2.591884e-10, -5.615886e-11, -1.728728e-11, 
    -2.432721e-13, -7.762679e-12, -4.146905e-12, 7.265299e-13, 3.394018e-11, 
    7.148282e-12, 2.300182e-11, 4.338774e-11, 3.150391e-11, 1.960754e-10, 
    4.435081e-10, -1.21757e-10, 5.005751e-11, -7.549583e-11, -2.326341e-10, 
    -1.150109e-10, 1.140166e-10, -3.723266e-11, 1.411249e-11, 2.593941e-10, 
    -1.599123e-10, 1.560663e-12, -2.362555e-13, 5.160306e-10, -5.049294e-14, 
    -1.694098e-11, 3.413336e-11, 2.073042e-11, -8.375661e-13, 1.385609e-10, 
    6.397127e-11, 1.250999e-12, 2.663314e-12, 2.146772e-12, 2.211842e-13, 
    4.308831e-11, -7.949841e-11, -6.620349e-12, 4.776135e-12, 3.470557e-13, 
    2.779998e-13, 2.495286e-10, -9.160672e-13, -1.609424e-11, -7.840673e-12, 
    -3.882072e-11, 6.757639e-11, -1.65572e-11, -5.821166e-12, -8.917711e-12, 
    1.025525e-09, -1.105671e-11, -4.657259e-10, -1.564058e-10, 6.961343e-11, 
    -9.039991e-11, 1.245437e-10, 1.393345e-10, -6.499534e-11, -9.010526e-12, 
    3.885781e-14, 5.884182e-15, -2.084055e-11, -3.415279e-12, 5.737211e-11, 
    -7.615464e-12, 5.007506e-12, 3.624434e-12, -1.096414e-10, -1.289613e-11, 
    -3.288718e-10, 1.108764e-10, 5.025691e-11, 1.028191e-12, -1.948885e-12, 
    -3.051537e-11, 8.98881e-13, 1.875389e-12, -1.755684e-11, -3.194178e-11, 
    -1.35806e-11, -8.548939e-12, 1.681388e-11, -6.009615e-11, -2.084866e-12, 
    4.924128e-11, 4.003362e-11, -8.418266e-14, 7.255863e-13, 9.568124e-12, 
    4.603451e-11, -5.262235e-12, -2.070322e-11, -3.051115e-12, 1.133249e-11, 
    -1.810929e-11, -1.090439e-11, -2.74869e-12, 3.63245e-11, 1.143996e-11, 
    4.098944e-14, 5.400125e-13, 3.936157e-13, 1.152856e-12, 5.738987e-11,
  -8.138823e-12, 3.555911e-11, -5.46132e-11, -1.469935e-12, 9.438894e-11, 
    7.636558e-11, -6.797141e-11, -3.383676e-10, -7.750911e-11, -4.554623e-11, 
    1.204339e-10, -9.722889e-12, 2.377591e-10, -9.55378e-11, 3.831024e-11, 
    -6.273204e-13, -7.642508e-12, -4.381384e-12, 1.657008e-11, 4.314638e-11, 
    2.612577e-12, 4.637002e-11, -7.323298e-11, -1.319984e-10, 5.149436e-11, 
    9.31033e-11, 1.83678e-10, 6.519896e-11, -2.240665e-10, -2.157901e-10, 
    -2.665757e-10, 2.324287e-10, 4.694378e-11, 7.874812e-11, 3.531291e-10, 
    -5.263585e-10, 3.976197e-12, -2.043921e-13, 4.339658e-10, 1.06799e-12, 
    -5.776144e-11, 3.458878e-11, 1.489653e-11, -1.677485e-12, 3.829883e-10, 
    3.863532e-11, 6.232348e-12, 9.950818e-12, -3.636025e-12, -1.216194e-12, 
    5.730472e-11, -7.238787e-11, -1.751181e-11, -3.739142e-12, 1.019651e-12, 
    2.033929e-13, 3.181078e-10, -2.675194e-13, -3.481855e-11, -3.995604e-11, 
    -6.076117e-11, 1.154326e-10, -1.972866e-11, -9.827072e-12, -7.953194e-12, 
    -2.310374e-11, -3.731593e-11, -2.543716e-10, -2.314966e-10, 8.271961e-11, 
    -1.813061e-10, 6.241319e-11, 3.66525e-10, -1.338085e-11, -1.765969e-11, 
    7.904788e-14, 2.892131e-14, -3.708334e-11, -3.023692e-12, 7.780532e-11, 
    -6.394441e-12, -7.4867e-12, 2.366551e-12, -2.278409e-10, -6.327974e-10, 
    1.771157e-10, 9.048762e-12, 6.249889e-11, 6.073288e-12, -2.876144e-12, 
    7.314149e-13, 3.071277e-11, 1.493472e-12, 6.939516e-12, -4.647882e-11, 
    -1.035563e-11, 7.818457e-12, -2.769829e-11, -3.787015e-11, -1.75957e-12, 
    1.109504e-10, 8.988776e-11, -3.037015e-13, 1.177503e-12, 4.662271e-11, 
    1.054112e-10, 3.983214e-11, 3.809975e-11, 8.792078e-12, 2.341238e-11, 
    -1.742517e-11, -1.342926e-11, 8.504752e-12, 4.986767e-11, -5.443646e-12, 
    6.155077e-14, 1.273148e-12, -1.020295e-13, 1.013606e-12, 2.20536e-10,
  -2.067191e-11, -1.730127e-11, -5.971668e-12, 1.422555e-10, 7.382939e-11, 
    -3.083356e-11, -2.90723e-11, -4.238383e-10, -1.399427e-10, -4.149263e-10, 
    -1.204286e-10, 1.649876e-10, 3.437495e-10, -1.257141e-10, 1.456262e-10, 
    6.872725e-13, -3.819789e-12, 1.449063e-12, 2.929834e-11, 4.063727e-11, 
    -8.699708e-13, 7.987166e-11, -1.381433e-10, -4.895555e-10, 1.328888e-10, 
    5.497958e-11, 3.570304e-10, 3.835376e-11, -4.027467e-10, -2.677507e-10, 
    -1.397624e-10, -3.838219e-11, 8.784307e-11, 4.606115e-10, 3.698521e-10, 
    -3.463652e-10, 8.995293e-12, -1.858513e-13, 2.297944e-10, 6.005152e-12, 
    -1.514091e-10, 3.658185e-11, 4.186651e-12, -2.109035e-12, 1.128337e-10, 
    -1.344245e-10, 1.2923e-11, 2.74738e-11, -1.775424e-11, -4.442446e-12, 
    5.999734e-11, -1.574638e-10, -2.803544e-11, -2.535705e-11, 1.279066e-12, 
    -3.761436e-13, -2.435963e-11, 7.522871e-13, -8.949001e-11, -1.047671e-10, 
    -7.837064e-11, 1.299347e-10, 1.182743e-11, -7.190604e-12, 2.495159e-12, 
    -1.137725e-10, -4.090017e-11, -3.389009e-10, -6.658007e-11, 6.558887e-11, 
    -2.235923e-10, 1.247891e-13, 2.150657e-10, 9.924639e-11, -3.499841e-11, 
    -3.370637e-13, 7.671641e-14, -2.978839e-11, 3.23257e-12, 9.25815e-11, 
    -7.004175e-12, -7.880785e-12, 1.718625e-13, -3.083094e-10, -3.05671e-11, 
    8.577019e-10, -2.828537e-11, 7.899326e-11, 1.650641e-11, 1.396527e-11, 
    3.309308e-11, 1.777378e-11, 1.826095e-12, 1.33122e-11, -5.541656e-11, 
    6.746337e-12, 1.44273e-11, -1.136686e-10, -8.640644e-12, 2.096901e-12, 
    1.324589e-10, 2.269863e-10, -4.815592e-13, 1.462441e-12, 3.739009e-11, 
    1.42113e-11, -1.203735e-10, -6.316236e-11, -8.01581e-13, 2.504885e-11, 
    -1.002887e-11, -1.345546e-11, 2.538014e-11, 4.548228e-11, -4.118972e-11, 
    1.000977e-13, 1.866174e-12, 5.380696e-13, -6.139533e-13, 2.875455e-10,
  -1.29301e-11, -2.726352e-11, 1.173888e-10, 1.26029e-10, -9.983658e-11, 
    8.514078e-12, 2.30612e-10, -3.526122e-10, -1.747935e-10, -7.992362e-10, 
    -4.144436e-10, 2.488498e-10, 9.092691e-10, -1.497202e-10, 1.596181e-10, 
    3.699618e-12, 2.843059e-12, 4.851231e-12, 3.091549e-11, 5.232792e-11, 
    -2.879474e-12, 8.719248e-11, -8.173018e-12, -6.16307e-10, 5.710188e-10, 
    5.561507e-10, 3.862297e-10, -3.071499e-11, -6.970389e-10, -2.988596e-10, 
    2.89706e-11, -2.120828e-10, -1.536549e-12, -3.098553e-10, 1.823306e-10, 
    -6.6788e-10, 1.351292e-11, -1.039169e-13, 2.954792e-10, 1.425455e-11, 
    -3.259892e-10, 2.067679e-11, -3.842704e-12, -8.056361e-12, 5.818226e-10, 
    -1.353833e-10, 1.778222e-11, 7.452261e-11, -3.726406e-11, -8.472223e-12, 
    3.214162e-11, -3.001883e-10, -3.856311e-11, -3.485283e-11, 1.434408e-14, 
    -5.719869e-13, -5.938041e-10, 1.417355e-12, -1.854016e-10, -2.517391e-10, 
    -9.570478e-11, 1.107008e-10, 1.185168e-10, 3.261391e-13, 1.246185e-11, 
    -2.078338e-10, 4.201617e-10, -7.149019e-10, -2.176783e-10, -3.430145e-12, 
    -2.74829e-10, -1.385114e-10, 3.743672e-11, 1.64615e-11, -5.444001e-11, 
    -4.263256e-13, 1.751932e-13, -9.462653e-12, 1.424256e-11, 1.240092e-10, 
    -1.490363e-11, -1.996581e-12, -3.17435e-12, -3.958984e-10, 1.797709e-10, 
    1.206061e-09, -8.403411e-11, 9.560353e-11, 4.517328e-11, 7.144862e-11, 
    -3.467271e-11, -1.46963e-10, 3.28626e-12, 4.451728e-12, -1.533884e-11, 
    3.450662e-11, 8.66045e-12, -1.820055e-11, 6.608047e-12, 5.326584e-12, 
    4.895817e-11, 4.083823e-10, -9.936496e-14, 3.777312e-12, -1.1166e-10, 
    -4.595968e-11, -1.576872e-10, -3.125074e-10, 3.902301e-11, 2.686384e-11, 
    3.964828e-12, -1.075939e-11, 2.692779e-11, 4.13749e-11, -7.000267e-11, 
    7.458922e-13, 1.933342e-12, 1.97703e-12, -4.146461e-12, 2.687308e-10,
  5.771383e-12, 8.639667e-11, 2.741327e-10, 1.402949e-10, -1.356621e-10, 
    -7.302425e-11, 4.762342e-10, -1.683489e-10, -2.102976e-10, -9.683863e-10, 
    3.03082e-11, 7.65958e-10, 2.077902e-09, -1.968115e-10, -2.749267e-11, 
    7.358736e-12, 1.64512e-11, 3.292477e-12, 1.881206e-11, 8.045475e-11, 
    -2.515321e-12, 6.311218e-11, -1.235456e-11, -1.082116e-09, 8.385541e-10, 
    1.043613e-09, 2.715357e-10, -4.493117e-10, -9.38476e-10, -2.015383e-10, 
    9.083756e-11, -7.825758e-10, -4.967973e-10, -7.300809e-10, 2.551381e-11, 
    -1.280878e-09, 5.678125e-12, 2.477796e-12, 4.762857e-10, 2.098677e-11, 
    -6.564534e-10, -3.015366e-11, -1.535794e-11, -1.684328e-11, 7.966143e-10, 
    -4.139444e-10, 1.956302e-11, 2.018212e-10, -6.957599e-11, -1.046996e-11, 
    2.980061e-11, -2.886029e-10, -5.430589e-11, -3.046843e-11, 6.77427e-12, 
    -3.907985e-13, -1.023444e-09, -4.91518e-13, -2.529351e-10, -2.914373e-10, 
    -1.174119e-10, 5.939071e-11, 2.599947e-10, 2.03606e-12, 1.259934e-11, 
    -8.48619e-11, -3.078569e-10, -1.01765e-09, -6.430234e-11, -1.603855e-10, 
    -5.998384e-10, -3.504113e-10, 4.72129e-10, -4.098393e-10, -5.655298e-11, 
    -3.462119e-12, 4.094503e-13, 5.221601e-12, 2.545058e-11, 2.007354e-10, 
    -2.340439e-11, 7.320069e-11, -4.97824e-12, -7.746941e-10, 3.459881e-10, 
    9.555947e-10, -3.513314e-10, 1.016645e-10, 1.084566e-10, 1.712355e-10, 
    -1.433751e-10, -1.785697e-10, 4.643841e-12, -9.633769e-11, 1.503118e-10, 
    5.231264e-11, -1.951719e-11, 2.181064e-10, 3.066525e-11, 9.745804e-12, 
    -1.237819e-10, 4.454394e-10, 1.94289e-12, 1.44732e-11, -3.818581e-10, 
    -1.725233e-10, 2.302603e-10, -2.492726e-10, 5.662955e-10, 8.199308e-11, 
    2.147971e-11, -9.84457e-12, 2.460077e-11, 1.028493e-10, -8.030909e-11, 
    2.831158e-12, 1.70397e-12, 4.116707e-12, -6.687095e-12, 2.179128e-10,
  -2.76863e-11, 4.072582e-10, 3.830749e-10, 3.293827e-10, 1.158149e-10, 
    -1.954312e-10, 2.944915e-10, 5.247713e-11, -3.34623e-10, -1.008608e-09, 
    7.094307e-10, 1.518856e-10, 1.023523e-09, -3.226432e-10, -9.781687e-11, 
    9.102052e-13, 3.232437e-11, 4.760636e-12, 3.622436e-12, 1.008154e-10, 
    4.618528e-13, 5.980283e-11, -6.859224e-11, -2.246399e-09, 5.806875e-10, 
    1.447493e-09, -4.709122e-11, -1.199645e-10, -1.930545e-10, -5.862368e-10, 
    -2.323297e-10, -5.4834e-10, -1.244917e-09, -2.029498e-09, 1.43352e-11, 
    -1.951779e-09, -3.174456e-11, 9.222845e-12, 3.713687e-10, 3.627143e-11, 
    -2.166985e-10, -8.167689e-11, -3.750245e-11, -2.906747e-11, 7.587033e-10, 
    -1.075538e-09, 3.531397e-11, 5.115632e-10, -1.135462e-10, -1.905542e-11, 
    4.51581e-10, -4.838796e-12, -1.018215e-10, -3.966889e-11, 3.809628e-11, 
    -2.73559e-13, -1.361599e-09, -8.199663e-13, -1.947527e-10, 8.756547e-10, 
    -1.705978e-10, 1.753975e-11, 2.095852e-10, -4.730083e-12, 6.570388e-12, 
    8.179413e-10, 2.070035e-09, -1.125073e-09, 4.548895e-10, -3.319442e-10, 
    -1.476359e-09, -4.627481e-10, 7.167387e-10, -7.790462e-10, -2.82423e-11, 
    -7.691625e-12, 5.511147e-13, 1.597744e-11, 4.08634e-11, 3.593215e-10, 
    -2.503597e-11, 2.354935e-10, -8.608225e-12, -9.571721e-10, -4.390444e-10, 
    4.971383e-10, -5.236913e-10, 9.627854e-11, 1.984406e-10, 2.622578e-10, 
    -2.251497e-10, -1.954383e-10, 4.6807e-12, -2.683468e-10, 5.894734e-10, 
    3.307328e-11, -6.439507e-11, 3.314113e-10, 3.173639e-11, 2.402913e-11, 
    -2.05997e-10, 3.654883e-10, 4.964251e-12, 3.996936e-11, -6.798473e-10, 
    -6.006715e-10, 1.414548e-10, 4.697895e-10, 1.35471e-09, 3.261711e-10, 
    4.200373e-11, 2.613731e-11, -1.666223e-12, 1.469083e-10, -6.20517e-11, 
    6.727774e-12, 2.249312e-12, 5.983103e-12, -8.010481e-12, 1.647145e-10,
  -2.792113e-10, 5.301253e-10, 4.658922e-10, 5.403145e-10, 2.937206e-10, 
    3.625722e-10, -4.469136e-10, 6.509318e-10, -5.72296e-10, -1.329379e-09, 
    8.980727e-10, -6.487362e-10, -4.212904e-09, -5.074376e-10, -2.527081e-10, 
    -1.284839e-10, 3.032525e-11, 1.32232e-11, 2.606804e-11, 9.441337e-11, 
    7.819523e-12, 7.222312e-11, 1.967138e-11, -1.668649e-09, 2.70223e-10, 
    2.818613e-09, -4.626379e-10, -6.275158e-11, -4.652385e-10, -1.064638e-09, 
    -9.295142e-10, -1.935696e-10, -1.995527e-09, -2.676185e-09, 2.859935e-12, 
    -1.810783e-10, -6.776943e-11, 1.727862e-11, -7.464855e-10, 1.721233e-10, 
    1.769202e-10, -6.141576e-11, -3.842615e-11, -5.071343e-11, 7.83853e-10, 
    -1.628482e-09, 1.012062e-10, 1.052223e-09, -1.462119e-10, -4.750511e-11, 
    1.172326e-09, -1.567777e-10, -2.151147e-10, -8.538592e-12, 7.595258e-11, 
    -8.277823e-13, -5.748468e-10, 7.372591e-12, -5.3776e-11, 2.827836e-10, 
    -2.642189e-10, -2.76934e-11, -7.54703e-11, -1.844214e-11, -3.716849e-12, 
    3.335412e-09, 1.12988e-09, -1.65355e-09, -1.794614e-09, -2.794813e-10, 
    -2.389942e-09, -5.290453e-10, 9.929799e-10, -1.247567e-09, -1.155556e-11, 
    -3.719691e-12, 1.254996e-12, 3.907452e-11, 6.14607e-11, 3.573781e-10, 
    -1.95044e-12, 2.910907e-10, -1.502443e-11, -6.667555e-10, -4.456812e-09, 
    -1.337224e-09, -6.516139e-10, 8.101964e-11, 2.483878e-10, 3.06315e-10, 
    -3.908589e-10, -3.534829e-10, 1.755041e-12, -3.319116e-10, 1.96739e-09, 
    -1.487805e-11, -1.050701e-10, 5.948309e-11, 7.300827e-12, 5.397922e-11, 
    -1.443574e-10, 9.84941e-11, -4.458656e-13, 7.703127e-11, -7.747794e-10, 
    -1.265544e-09, -8.456063e-10, 7.046985e-10, 3.833911e-10, 6.716867e-10, 
    6.99778e-11, 4.215295e-11, 3.776535e-12, 1.21414e-10, -7.016965e-11, 
    1.200959e-11, 3.61311e-12, 5.717427e-12, -8.502976e-12, 9.780265e-11,
  -4.616219e-10, 7.567458e-10, 2.048896e-09, -5.834515e-10, -8.826468e-10, 
    5.988205e-10, -2.376872e-10, 1.190333e-09, -9.67102e-10, -8.244534e-10, 
    3.194209e-10, -1.833307e-10, -1.839577e-09, -6.533689e-10, -4.133902e-10, 
    -7.501406e-10, -5.952145e-11, 4.477485e-11, 8.579448e-11, 9.712053e-11, 
    2.969003e-11, 2.007283e-12, 7.44258e-11, 5.351417e-10, 9.140777e-11, 
    5.180613e-09, 1.069555e-09, -2.556202e-09, -7.795045e-10, 1.739071e-09, 
    -5.813089e-09, -5.895622e-10, -2.470568e-09, 2.502876e-09, -3.899103e-11, 
    -1.850079e-09, -2.729124e-11, 2.098766e-11, -1.420442e-09, 6.589154e-10, 
    9.519639e-11, 3.865708e-11, 1.966782e-11, -1.552576e-10, 9.157937e-10, 
    -1.688175e-09, 2.010161e-10, 1.459188e-09, -3.100176e-10, -5.221956e-11, 
    9.859953e-10, -2.477343e-10, -3.514536e-10, 1.643777e-10, 7.721361e-11, 
    -2.312817e-12, -1.695991e-09, 2.297966e-11, -2.609468e-11, 2.176037e-12, 
    -3.564899e-10, -1.279368e-10, -1.152891e-10, -2.140936e-11, 
    -1.723137e-11, 7.579178e-09, -4.569753e-09, -4.733348e-09, -2.39184e-09, 
    -1.677698e-10, -2.173362e-09, 3.411351e-10, 5.194387e-10, -2.007962e-09, 
    7.235243e-11, 9.553247e-12, 3.712586e-12, 8.509105e-11, 7.505463e-11, 
    -2.180904e-10, 5.901413e-11, 4.773085e-10, -2.576073e-11, 4.947829e-10, 
    -4.114138e-09, -2.232493e-09, -7.160814e-10, 5.259793e-11, 3.141452e-10, 
    2.415881e-10, -9.303953e-10, -8.524374e-10, -6.110668e-12, -4.504635e-10, 
    1.712625e-09, -9.901484e-11, -1.384386e-10, -3.14099e-10, -9.972467e-12, 
    1.145857e-10, -6.878587e-10, -2.61239e-10, -1.497824e-11, 1.172564e-10, 
    -8.010339e-10, -1.676806e-09, -1.437709e-09, 3.096297e-10, -4.182606e-09, 
    1.124494e-09, 3.911538e-12, -8.71232e-11, 5.228529e-11, 1.109335e-10, 
    -1.413945e-10, 2.230891e-11, 8.121503e-12, 4.19309e-12, -8.871126e-12, 
    1.829292e-11,
  -5.975593e-10, 4.260734e-09, 4.051451e-09, -1.767994e-09, -4.762263e-09, 
    -3.597343e-09, 1.455042e-09, 6.522711e-10, 4.046896e-10, 6.900009e-10, 
    8.471801e-11, 1.178513e-09, -1.167969e-09, -7.189342e-10, -6.926584e-10, 
    -1.398752e-09, -3.975586e-10, 6.296119e-11, 1.058531e-10, 2.357794e-10, 
    7.371881e-11, -8.981971e-11, 1.21112e-10, 2.141199e-09, -4.041354e-10, 
    4.681461e-09, 2.541888e-09, -5.808197e-09, -9.454268e-10, 1.947889e-09, 
    -1.567464e-09, -6.263434e-11, -1.015458e-09, 1.445123e-09, 4.546763e-11, 
    -3.010591e-09, 5.992717e-11, 2.927436e-11, -3.210637e-09, 1.473982e-09, 
    -5.068913e-10, 1.50564e-11, 9.667644e-11, -4.648875e-10, 2.161038e-09, 
    -1.032184e-09, 2.393747e-10, 1.42288e-09, -8.973714e-10, -4.143974e-11, 
    6.355432e-10, -8.244356e-10, -2.304802e-10, 3.754778e-10, 9.915411e-11, 
    -2.209788e-12, 1.471754e-09, 4.120864e-11, -1.681514e-10, 1.416804e-10, 
    -3.509726e-10, -1.924505e-10, -3.806377e-11, -3.488339e-11, 
    -2.072653e-11, 1.382605e-08, 6.72479e-10, 2.326722e-09, -3.06455e-09, 
    -5.163869e-10, 4.587193e-10, 1.777927e-09, 1.205294e-10, -2.086288e-09, 
    1.47152e-10, 3.463896e-11, 1.260858e-11, 1.673008e-10, 3.330172e-11, 
    1.477289e-10, 2.328164e-10, 9.843277e-10, -2.037837e-11, 2.014183e-09, 
    -2.489436e-09, 5.576126e-10, 9.645618e-11, 3.056044e-11, 6.134528e-10, 
    -1.861622e-11, -2.092982e-09, -1.250324e-09, -1.4726e-11, -6.725188e-10, 
    2.576762e-09, -1.494897e-10, -1.101355e-10, -2.947971e-10, -2.045653e-11, 
    1.575685e-10, -1.636487e-09, -6.811796e-10, -2.902656e-11, 1.60493e-10, 
    -1.276867e-09, -1.860862e-09, -1.692818e-09, -3.497362e-10, 
    -3.985399e-09, 2.111172e-09, 5.122303e-11, -3.196092e-10, 1.152145e-10, 
    -4.357403e-10, -2.859863e-10, 3.258123e-11, 1.968203e-11, 6.785239e-12, 
    -1.28626e-11, -4.17586e-11,
  -6.309264e-10, 6.371302e-09, 5.91605e-10, -3.255352e-10, 1.823629e-09, 
    -1.251947e-08, 1.283844e-09, -7.525713e-10, 1.534268e-09, 1.95076e-09, 
    7.597478e-10, 3.810335e-09, -7.126744e-12, -7.674359e-10, -9.266259e-10, 
    -1.409784e-09, -1.798388e-09, 6.321699e-11, -4.263256e-13, 3.452456e-10, 
    1.105676e-10, -1.421299e-10, -1.144684e-11, 1.55061e-09, 8.931522e-12, 
    -2.175042e-10, 4.554245e-09, -8.361717e-09, -3.987211e-10, 3.037322e-09, 
    -8.738475e-09, 8.525447e-10, 1.75681e-09, 2.034717e-09, 2.567688e-10, 
    -9.863776e-09, 2.7201e-11, 2.770406e-11, -6.339228e-09, 2.308458e-09, 
    -1.262099e-09, -2.620695e-10, 1.259792e-10, -2.626255e-10, 3.252559e-09, 
    -9.539391e-10, 1.520775e-10, 1.213287e-09, -1.694978e-09, -5.235101e-11, 
    1.060503e-09, -1.226589e-09, 5.137551e-10, 4.656002e-10, 2.545136e-10, 
    2.053469e-12, 5.270302e-09, 5.801013e-11, -4.502269e-10, 5.257839e-10, 
    -2.290435e-10, -1.981206e-10, -1.744382e-11, -4.206456e-10, 
    -4.144312e-11, 1.107887e-08, 1.384542e-09, 3.2909e-09, -4.946422e-09, 
    -1.615142e-09, 6.951453e-10, 3.001624e-09, 3.203482e-10, -2.402309e-09, 
    -9.338365e-10, 1.003642e-10, 1.86624e-11, 3.554277e-10, -6.825189e-11, 
    6.727205e-10, 5.600995e-10, 9.691185e-10, 4.147438e-11, 4.178254e-09, 
    1.231292e-09, 6.586234e-10, 1.826557e-09, 3.530687e-11, 2.530229e-10, 
    4.973302e-10, -3.316011e-09, -2.819761e-10, -2.368949e-11, -1.720061e-09, 
    2.433843e-09, -9.982699e-11, 7.725162e-11, 6.741701e-10, -1.062617e-10, 
    2.430639e-10, -1.701231e-09, -9.25068e-10, -3.161205e-11, 2.019149e-10, 
    -2.849042e-09, -1.354401e-09, -2.152682e-09, 7.969234e-10, 2.036593e-09, 
    3.105306e-09, 2.342304e-10, -4.972591e-10, 1.474021e-10, -1.080018e-09, 
    -4.641194e-10, 4.187228e-11, 3.727862e-11, 2.295497e-11, -3.964296e-11, 
    -2.884093e-11,
  6.839613e-10, 8.100749e-09, -6.82909e-09, -9.657484e-10, -5.341924e-09, 
    -5.003507e-09, -5.436881e-09, 9.110224e-10, 1.49867e-09, 3.443056e-09, 
    1.155335e-09, 2.759826e-09, -6.271321e-10, -9.617125e-10, -1.369138e-09, 
    -9.558661e-10, -2.405169e-09, 2.012612e-10, -1.869793e-11, 4.481748e-10, 
    2.770193e-10, -1.497042e-10, -1.09516e-10, 2.202931e-09, 3.252225e-10, 
    -3.426528e-09, 6.36367e-09, -9.762296e-09, 2.327532e-09, 6.23006e-09, 
    -1.488176e-08, -2.251262e-09, 2.428372e-09, 5.08728e-09, 5.45576e-10, 
    -2.25517e-08, -3.357641e-10, 3.567635e-11, -9.306014e-09, 3.165023e-09, 
    -2.59284e-09, -5.889049e-10, -2.938378e-10, -2.186473e-10, 1.674714e-09, 
    -1.379824e-09, 7.769785e-11, 1.090363e-09, -2.104396e-09, 1.510614e-11, 
    1.244839e-09, -1.33074e-09, 4.186873e-10, 4.050818e-10, 5.462432e-10, 
    1.541878e-12, 3.091905e-09, 8.526371e-11, -8.130754e-10, -1.891756e-09, 
    -3.212293e-10, -2.518803e-10, 1.50564e-11, -1.254718e-09, 3.7587e-10, 
    1.599815e-08, -7.985435e-10, 2.320483e-09, 3.338009e-09, -2.302421e-09, 
    -1.010626e-09, 1.497874e-09, 4.615615e-10, -1.348788e-09, -2.215548e-09, 
    1.667146e-10, -8.675727e-12, 6.8529e-10, -1.112035e-10, -2.052118e-10, 
    1.117662e-09, -2.527328e-11, 1.593534e-10, 7.534872e-09, 5.724921e-09, 
    -7.228849e-10, 2.88005e-09, 8.804335e-11, 2.437983e-10, 1.333923e-09, 
    -3.754344e-09, 4.028593e-10, -2.656719e-11, -8.320298e-09, 7.235457e-11, 
    -9.521983e-11, 3.294517e-10, 1.822279e-09, -2.92836e-10, 2.89036e-10, 
    -5.154916e-10, -6.374457e-10, -2.640022e-11, 2.002309e-10, -1.77247e-09, 
    1.946816e-10, -2.003084e-09, -2.208147e-09, -8.527437e-10, 4.132566e-09, 
    4.351861e-10, -5.65457e-10, 3.68054e-10, -2.213177e-09, -6.654162e-10, 
    6.592842e-11, 6.841105e-11, 5.853984e-11, -1.11255e-10, -2.38245e-11,
  3.862063e-09, 6.489792e-09, 2.874465e-09, 2.273516e-09, -7.983587e-10, 
    -4.281695e-09, -1.571981e-08, 4.746774e-09, -5.799947e-10, 3.705004e-09, 
    2.899704e-09, 4.830625e-10, -5.649312e-10, -2.63114e-11, -2.076909e-09, 
    -6.135892e-10, -2.915284e-09, -7.62391e-10, 2.071943e-10, 8.425687e-10, 
    2.674838e-10, -1.377245e-10, -9.901413e-11, 1.665036e-09, -6.579839e-10, 
    -1.139277e-09, 6.604871e-09, -2.021149e-08, 3.030927e-09, 1.189188e-08, 
    -1.2723e-08, -7.169199e-09, -2.274803e-10, 6.656315e-09, 6.325891e-10, 
    -2.832578e-08, -6.635261e-10, 7.640111e-11, 3.233943e-09, 4.34461e-09, 
    -5.590515e-09, -9.166783e-10, -5.349392e-10, -2.935825e-10, 
    -3.383569e-09, -1.53198e-09, 8.950707e-11, 1.113321e-09, -2.305113e-09, 
    4.432117e-10, 2.218524e-09, -7.479954e-10, 3.481104e-10, 4.960512e-10, 
    8.570673e-10, -2.616929e-11, 3.588596e-10, 1.050509e-10, -6.331831e-10, 
    -1.37814e-09, -6.244747e-10, -4.390799e-10, 2.575362e-10, -6.219281e-10, 
    -1.613311e-09, 1.805297e-08, -4.036757e-09, 3.83757e-10, 1.203524e-09, 
    -2.413252e-09, 7.194743e-10, -4.176307e-09, 1.346976e-10, 2.74742e-09, 
    -1.209273e-10, 1.440768e-10, -5.965362e-11, 1.196156e-09, -1.714774e-10, 
    -1.463341e-09, 1.568246e-09, -1.586159e-10, 2.870948e-10, 1.024689e-08, 
    7.179104e-09, 2.834355e-11, 2.491085e-09, 2.254481e-10, 8.649046e-10, 
    2.129319e-09, -4.918228e-09, 6.947665e-12, -5.896794e-11, -1.935511e-08, 
    -1.009987e-09, -9.815011e-11, 4.831264e-11, 4.193126e-10, -5.747367e-10, 
    2.577295e-10, 4.93749e-10, 4.736638e-10, -1.885958e-11, 1.082388e-10, 
    9.200818e-11, 4.872405e-10, -7.785488e-10, -2.272081e-09, -1.507196e-09, 
    4.702947e-09, 3.009362e-10, -3.759553e-10, 7.862937e-10, -2.448949e-09, 
    -6.504237e-10, 7.342038e-11, 1.421263e-10, 8.995205e-11, -1.542251e-10, 
    -1.058922e-10,
  7.843994e-09, 5.14521e-09, 7.344312e-09, 9.627854e-10, 1.431232e-09, 
    2.296929e-09, -1.403458e-08, 4.296993e-09, 2.492584e-10, 2.578588e-09, 
    3.999816e-09, 1.703597e-09, -6.481855e-10, 2.024194e-09, 1.656161e-09, 
    -1.050924e-09, -5.339058e-09, -2.103477e-09, -1.067377e-10, 8.819825e-10, 
    2.875709e-10, 1.600426e-10, -1.138005e-10, 6.474465e-10, -1.632941e-09, 
    2.729678e-09, 5.925244e-09, -5.71541e-08, 1.102367e-08, 3.496942e-08, 
    -8.293455e-09, -4.827768e-09, -5.90191e-09, 7.704358e-09, 3.8537e-10, 
    -3.350377e-08, -9.590394e-10, 9.289991e-11, 1.810108e-08, 6.435357e-09, 
    -9.612575e-09, -1.50493e-09, -2.812754e-10, -5.066179e-10, -2.02985e-09, 
    -4.945349e-09, 1.026308e-10, 2.000242e-09, -2.623665e-09, 6.038015e-10, 
    2.768044e-09, -3.736034e-10, 3.101945e-10, 7.15886e-10, 1.175698e-09, 
    -7.463541e-11, -3.69937e-10, 1.827772e-10, -7.85056e-10, 5.66094e-09, 
    -6.722303e-10, -4.647802e-10, 6.123457e-10, -1.261867e-10, -6.996021e-09, 
    1.565951e-08, -4.962033e-09, 4.604885e-10, 5.405241e-10, -4.219999e-09, 
    3.162285e-09, -1.288467e-08, -6.386358e-10, 3.824994e-10, 6.152223e-09, 
    4.3201e-12, -1.256026e-10, 2.111385e-09, -2.34872e-10, 2.042952e-09, 
    2.101459e-09, 2.834512e-10, 4.384475e-10, 8.88474e-09, 4.2115e-09, 
    1.484352e-09, 9.66196e-10, 5.306049e-10, 1.394215e-09, 2.494062e-09, 
    9.869439e-10, -2.611898e-10, -1.195488e-10, -2.902535e-08, -1.966214e-10, 
    -9.008545e-11, -2.500065e-09, -3.139661e-09, -8.486438e-10, 8.922711e-11, 
    1.542588e-09, 2.130754e-09, -3.72129e-11, -3.553069e-11, 3.779235e-10, 
    6.498055e-10, 1.945182e-09, 1.368761e-09, -8.058407e-10, 3.626042e-09, 
    2.957279e-10, -1.213607e-11, 1.526814e-09, -2.83444e-09, -4.174296e-10, 
    -2.297895e-11, 2.764544e-10, 1.235136e-10, -1.526868e-10, -2.84416e-10,
  1.032191e-08, 5.803713e-11, -3.942091e-10, 3.728985e-09, 4.149967e-09, 
    3.210062e-09, -2.544709e-09, -1.759872e-09, 3.92356e-09, 5.032916e-10, 
    2.526747e-09, 8.07006e-10, 6.039045e-10, 2.856382e-10, 5.203049e-09, 
    -2.090218e-09, -7.372409e-09, -2.664734e-09, -9.850254e-10, 4.087042e-11, 
    2.049148e-09, 1.0549e-09, -2.884804e-10, 2.032721e-10, 3.22467e-09, 
    2.645436e-09, 6.308539e-09, -6.105108e-08, 1.919699e-08, 4.275807e-08, 
    -1.452696e-08, -5.69861e-09, -8.096947e-09, 8.460745e-09, -1.887202e-11, 
    -3.652553e-08, -1.542946e-09, 7.68452e-11, 5.580034e-09, 9.42394e-09, 
    -1.289635e-08, -2.618322e-09, -6.252776e-12, -6.844223e-10, 
    -1.045925e-08, -5.855668e-09, 5.062475e-10, 3.955449e-09, -3.44005e-09, 
    2.32351e-10, 2.486487e-09, -8.402594e-10, 5.277796e-10, 8.179996e-10, 
    1.579952e-09, -7.372591e-11, -3.986372e-09, -5.11136e-10, -2.048205e-09, 
    1.169636e-08, 8.866436e-10, -9.885071e-11, -6.872369e-11, -3.229013e-09, 
    -1.0339e-08, 2.156554e-08, -6.945925e-09, 7.651693e-10, -3.13031e-09, 
    -1.388457e-09, 3.068635e-09, 9.05851e-09, -2.122931e-09, -2.987406e-09, 
    1.491907e-08, -1.902549e-10, -1.861622e-10, 3.307619e-09, -3.140926e-10, 
    6.70866e-09, 3.243997e-09, 1.750868e-09, 5.712195e-10, 5.665299e-09, 
    -9.811174e-11, 3.641219e-09, -2.008733e-09, 8.013785e-10, 1.542062e-09, 
    2.639069e-09, 9.530993e-09, -6.974233e-10, -4.968115e-11, -2.434476e-08, 
    -1.341789e-09, -4.329763e-11, -5.738138e-09, -7.836206e-09, 
    -1.207923e-09, -2.380034e-10, -8.634515e-11, 3.311531e-09, -9.566392e-11, 
    -1.152358e-10, -7.08269e-11, 7.270273e-10, 1.452008e-09, 2.25009e-09, 
    -5.279617e-10, 7.820802e-09, 3.458581e-09, 1.704734e-10, 1.198202e-09, 
    -4.548838e-09, -7.739231e-10, -8.193411e-11, 3.572396e-10, 9.794654e-11, 
    -1.339515e-10, -6.609753e-10,
  9.807366e-09, -8.97785e-10, -1.546539e-09, 9.803216e-10, 1.192177e-09, 
    4.067715e-10, 2.377078e-09, -1.258582e-08, 5.473453e-09, -5.588845e-10, 
    1.058822e-09, 6.894538e-10, 1.785395e-09, -6.426433e-09, 6.534322e-09, 
    1.949957e-10, -8.726289e-09, -2.273879e-09, -1.641304e-09, -5.905463e-10, 
    3.795265e-09, 9.012524e-10, 8.071765e-11, -1.051035e-10, -1.096339e-09, 
    2.880483e-09, 1.962184e-08, -4.061962e-08, 1.80853e-08, 7.34525e-09, 
    -7.926019e-09, -6.784546e-09, -9.75632e-09, 1.001047e-08, 5.82645e-10, 
    -2.727052e-08, -2.008073e-09, 1.035687e-10, -4.477909e-08, 1.307505e-08, 
    -1.347039e-08, -3.995467e-09, -5.381651e-11, -1.021129e-09, -1.38017e-08, 
    -2.175511e-09, 1.092502e-09, 6.988088e-09, -4.564413e-09, 3.61851e-10, 
    1.859064e-09, -2.017373e-10, 4.027525e-10, 9.047313e-10, 2.056139e-09, 
    1.094236e-11, -3.001333e-09, -2.942113e-09, -3.438328e-09, 9.865801e-09, 
    3.518721e-09, 3.87729e-10, -1.707974e-09, -8.727488e-09, -2.408445e-09, 
    1.587392e-08, -9.135761e-09, -3.547825e-09, -4.782862e-09, 1.281819e-10, 
    1.703938e-09, 3.266928e-08, -1.643002e-09, 4.334936e-09, 1.971705e-08, 
    -4.227445e-10, -1.65052e-10, 4.514334e-09, -4.143985e-10, 1.498938e-08, 
    5.094819e-09, 3.852021e-09, 7.366907e-10, -2.659021e-09, 7.867698e-10, 
    2.784077e-09, -4.280594e-09, 8.886332e-10, 1.682325e-09, 2.550991e-09, 
    9.385872e-09, 1.941316e-10, 5.104539e-10, -6.054909e-09, -2.062848e-10, 
    -1.697345e-11, -6.482844e-09, -1.535756e-08, -1.741228e-09, 
    -6.384767e-10, -7.192398e-10, 2.275488e-09, -1.153317e-10, -2.214726e-10, 
    -1.935916e-09, 7.271979e-10, 1.246576e-09, 7.469794e-10, -1.749868e-09, 
    1.149039e-08, 5.327422e-09, 1.321609e-10, -8.150209e-10, -7.102358e-09, 
    -2.968477e-09, -7.806306e-11, 3.530758e-10, 6.914647e-11, -1.122444e-10, 
    -8.530492e-10,
  6.782727e-09, -1.01295e-09, -1.219291e-10, 1.791705e-10, -4.369554e-10, 
    -7.163976e-10, 3.300897e-10, -1.657759e-08, 3.204207e-09, 2.944944e-09, 
    -1.995772e-10, 6.599521e-11, 1.110607e-09, -6.001301e-09, -1.151932e-09, 
    -2.601098e-09, -1.085976e-08, -1.041769e-09, -2.715048e-09, 
    -5.946958e-10, 5.796494e-09, -3.699938e-10, 8.673737e-10, 7.622702e-11, 
    -1.158583e-09, -1.946091e-09, 3.132561e-08, -6.957231e-08, 1.088631e-08, 
    -7.232359e-09, -3.583807e-09, -8.923905e-09, -1.389367e-08, 1.376492e-08, 
    3.262414e-09, -1.595618e-08, -2.603349e-09, 1.472316e-10, -8.052587e-08, 
    1.804022e-08, -7.571714e-09, -2.806928e-09, -2.123812e-10, -1.488235e-09, 
    -1.276283e-08, -5.97629e-09, -2.277517e-09, 1.125173e-08, -5.133995e-09, 
    4.114327e-10, 1.457181e-09, 1.453657e-09, -4.029115e-10, 1.107548e-09, 
    2.458857e-09, 1.220144e-10, -6.005507e-09, -8.039915e-09, -4.776916e-09, 
    4.624312e-09, -2.1912e-09, 5.414904e-10, -3.573064e-09, -8.245922e-09, 
    4.644892e-09, 1.425394e-08, -1.028366e-08, -1.210651e-08, 1.249987e-09, 
    3.713012e-10, 3.300897e-10, 2.644526e-08, -3.639684e-10, 6.996061e-09, 
    1.465214e-08, -6.269261e-10, -4.467893e-11, 4.77938e-09, -6.203706e-10, 
    2.555146e-08, 6.984692e-09, 7.222427e-09, 9.928556e-10, -3.639116e-09, 
    5.227719e-09, 1.046658e-09, -1.268631e-09, 1.028582e-09, 1.967967e-09, 
    1.985853e-09, 8.173913e-09, 1.879039e-09, 1.38354e-09, 7.509984e-10, 
    1.128114e-09, -1.075932e-09, -6.42201e-09, -1.524734e-08, -3.171351e-09, 
    -1.025626e-09, 4.255298e-10, 2.883489e-10, -1.309992e-10, -3.561453e-10, 
    -7.221047e-09, -2.790614e-09, 1.371291e-09, -2.357524e-09, 4.399681e-11, 
    1.358836e-08, 4.00729e-09, 5.358061e-10, -3.539299e-09, -8.934762e-09, 
    -3.013668e-09, -2.670504e-11, 2.43233e-10, 3.326583e-11, -1.001617e-10, 
    -3.509513e-10,
  3.05522e-09, -1.741284e-09, 3.350351e-10, -1.401759e-10, -1.489695e-09, 
    -3.718696e-10, -4.074991e-09, -6.557343e-09, -1.106287e-09, 4.386436e-09, 
    1.279091e-09, -9.105179e-10, -2.672266e-09, 1.261469e-09, -1.430828e-08, 
    -3.792127e-09, -1.519525e-08, 2.479396e-09, -4.861043e-09, -2.043521e-10, 
    8.790835e-09, 1.558874e-09, 4.633876e-10, 1.171998e-09, 3.74655e-10, 
    -2.256343e-09, 2.264505e-08, -4.061638e-08, -1.239329e-08, 1.67214e-08, 
    -1.383e-10, -1.11533e-08, -1.955971e-08, 1.636658e-08, 4.602555e-09, 
    -1.336718e-08, -2.21695e-09, 1.619966e-10, -6.468196e-08, 2.346063e-08, 
    1.321313e-09, 3.444882e-09, 2.080469e-11, -2.471267e-09, -2.980579e-08, 
    -1.569492e-08, -1.416413e-08, 1.758391e-08, -4.751598e-09, 4.652172e-10, 
    9.572503e-10, 1.386866e-09, 7.127397e-09, 9.878818e-10, 2.994374e-09, 
    1.866454e-10, -1.212328e-08, -1.748579e-08, -1.023578e-08, -9.49219e-09, 
    -1.353743e-08, 1.371291e-09, -3.224272e-09, -1.317892e-09, 4.86084e-09, 
    2.347298e-08, -2.324498e-09, -2.949145e-08, 4.694414e-09, 1.857813e-09, 
    2.529532e-10, 1.978833e-09, 3.029754e-11, 2.178695e-09, 6.92026e-09, 
    -6.522214e-10, -4.26752e-11, 3.897298e-09, -9.423743e-10, 2.902419e-08, 
    8.315169e-09, 1.270776e-08, 1.355318e-09, -3.636671e-09, 1.009056e-08, 
    5.418315e-10, 2.171248e-09, 9.530368e-10, 2.15081e-09, 2.712966e-09, 
    9.694077e-09, 5.488198e-09, 2.090388e-09, -7.162145e-09, 2.268166e-09, 
    -5.318907e-09, -7.502171e-09, 5.599361e-09, -5.633922e-09, -1.315777e-09, 
    -3.527703e-10, -2.360068e-10, -3.778347e-10, -3.175238e-10, 1.526928e-09, 
    2.085528e-09, 4.118647e-09, -4.067033e-09, 6.312462e-09, 1.179103e-08, 
    1.275737e-09, -1.772378e-10, -4.170715e-09, -1.152932e-08, -1.393119e-09, 
    4.127969e-11, -4.156675e-11, -2.246381e-11, -1.002896e-10, 4.914682e-10,
  7.531753e-10, -7.123617e-10, -5.944685e-10, -1.257376e-09, -2.052957e-09, 
    -1.570413e-09, -7.542042e-09, 4.684125e-09, -1.11973e-08, 7.632366e-10, 
    3.799755e-09, -1.359808e-09, -4.428387e-09, 3.295895e-09, -4.664003e-09, 
    -4.697239e-09, -1.775289e-08, 6.592046e-09, -9.165852e-09, -1.294325e-10, 
    1.051149e-08, -1.947228e-09, 1.211504e-09, 2.374122e-09, 1.622709e-09, 
    -6.660343e-10, -1.270223e-08, -2.861418e-08, -5.144955e-08, 2.235998e-08, 
    -5.811557e-09, -1.361821e-08, -2.363043e-08, 2.170924e-08, 3.295611e-09, 
    2.296076e-08, -1.00481e-09, 1.795897e-10, -4.986214e-08, 2.443648e-08, 
    1.12545e-08, 6.017046e-09, 9.316494e-10, -2.788331e-09, -4.634302e-08, 
    -1.964344e-08, -3.212435e-08, 2.666501e-08, -3.402806e-09, 3.975131e-10, 
    -4.395332e-09, -1.368903e-09, 1.086456e-08, 7.027552e-10, 3.887299e-09, 
    1.980709e-10, -2.063138e-08, -2.178947e-08, -1.8684e-08, -1.953465e-08, 
    -5.578841e-09, 2.197453e-09, -1.226283e-09, 6.953928e-09, 7.580753e-09, 
    2.667139e-08, 9.109442e-09, -2.98819e-08, 1.06175e-08, 5.152515e-09, 
    -5.390348e-09, -3.111552e-09, -8.907477e-09, -1.420858e-09, 3.687478e-09, 
    -6.05894e-10, 4.631318e-11, 3.488864e-09, -1.371775e-09, 1.883188e-08, 
    8.128637e-09, 2.159011e-08, 1.800316e-09, -8.390089e-11, 1.953936e-09, 
    -7.167387e-10, 4.367735e-09, 9.663381e-12, 1.324807e-11, 5.614368e-09, 
    1.16874e-08, 8.078302e-09, 2.361077e-09, -1.986923e-08, 1.436945e-09, 
    -1.037264e-08, -9.307416e-09, 2.27468e-08, -6.145513e-09, -1.458955e-09, 
    -1.287276e-09, -9.059207e-10, -8.489742e-10, -9.51772e-11, 1.241966e-08, 
    4.216417e-09, 2.695003e-09, 7.689209e-10, 8.228028e-09, 5.171216e-09, 
    -1.716899e-09, -1.285855e-09, -8.014922e-11, -1.725982e-08, 
    -7.158064e-09, 1.419664e-10, -5.641638e-10, -9.062973e-12, -1.050502e-10, 
    2.889976e-09,
  -2.9479e-10, 3.051355e-10, -6.540404e-10, -1.908006e-09, -1.148237e-09, 
    -3.275886e-09, -9.92236e-09, 9.286111e-09, -2.159857e-08, -7.825122e-09, 
    -5.210268e-10, -2.111562e-09, 7.319159e-10, 1.120952e-10, 6.686832e-09, 
    -5.206817e-09, -1.964494e-08, 9.037848e-09, -1.606328e-08, -1.307342e-09, 
    9.902749e-09, -2.137369e-09, 3.270657e-09, 2.09036e-09, 1.773287e-09, 
    3.685159e-10, -9.53533e-08, -2.397348e-08, -1.210917e-07, 2.933263e-08, 
    -8.561983e-09, -1.769081e-08, -2.330984e-08, 3.506835e-08, 1.014428e-09, 
    3.313056e-08, 2.07699e-09, 2.786962e-10, -4.473412e-08, 1.954741e-08, 
    2.247501e-08, 4.407298e-09, 2.224098e-09, -4.399453e-09, -4.208636e-08, 
    -1.83885e-08, -4.850122e-08, 4.024207e-08, -7.339964e-10, 2.644605e-10, 
    -7.283411e-09, -5.077368e-09, 3.115201e-08, 7.340076e-10, 5.276547e-09, 
    1.608953e-10, -3.471769e-08, -2.192915e-08, -2.932293e-08, 7.913314e-11, 
    7.938013e-09, 1.230831e-09, -1.609465e-09, 9.641508e-09, 8.62757e-09, 
    2.561467e-08, 1.221343e-08, 4.184545e-08, 1.057595e-08, 3.806349e-09, 
    -4.518762e-08, 3.413106e-09, 6.747484e-09, -3.094669e-09, 8.68418e-09, 
    -2.373213e-10, 3.24377e-10, 1.522324e-09, -2.174177e-09, 6.276082e-09, 
    8.818859e-09, 3.375499e-08, 2.328562e-09, 6.486403e-10, 3.56863e-10, 
    -2.213028e-09, 7.495601e-09, -1.940066e-10, 7.104147e-09, 1.162783e-08, 
    7.287326e-09, 4.165383e-09, 2.157407e-09, -6.959494e-09, 3.525429e-10, 
    -1.983657e-08, -1.325087e-08, 8.260258e-09, -8.752636e-09, -1.560215e-09, 
    -2.37128e-09, 3.639435e-10, -1.575771e-09, 1.387654e-10, 2.725301e-09, 
    -2.18165e-10, 9.003998e-11, 1.154717e-09, 3.89781e-09, 1.424155e-09, 
    -3.251728e-09, -6.293135e-10, 1.533465e-09, -2.162852e-08, -1.481629e-08, 
    2.593879e-10, -2.141363e-10, 7.535306e-12, -5.663381e-11, 5.286267e-09,
  -2.879858e-09, -2.268052e-11, 2.232241e-09, -1.033527e-09, -3.703917e-10, 
    -1.887884e-09, -9.817541e-09, 2.438071e-09, -2.076331e-08, -1.496028e-08, 
    -5.466291e-09, 4.874892e-10, 2.025956e-09, 1.64755e-09, 2.347792e-08, 
    -4.913386e-09, -2.162973e-08, 9.414777e-09, -2.429056e-08, -3.433627e-09, 
    1.137744e-08, 3.564821e-09, 7.95751e-10, 1.473438e-09, 1.0034e-09, 
    6.064624e-10, -6.295295e-09, -2.292808e-08, -1.611746e-07, 5.356134e-08, 
    -1.96755e-08, -1.333905e-08, -2.236663e-08, 4.715542e-08, 1.904425e-09, 
    4.4476e-08, 3.445319e-09, 5.457537e-10, -4.035519e-08, 5.732272e-09, 
    4.793979e-08, 4.032017e-09, 3.152977e-09, -1.197765e-08, -1.791955e-08, 
    -5.660593e-08, -5.85041e-08, 5.439001e-08, 1.833689e-09, 2.21128e-10, 
    -2.154543e-09, -2.96933e-09, 4.953596e-08, 1.328146e-09, 7.251306e-09, 
    8.242296e-12, -5.364672e-08, -1.111329e-08, -5.259191e-08, 3.466854e-08, 
    9.521727e-09, -7.083258e-10, -3.243542e-09, 7.854874e-09, 8.547874e-09, 
    2.259964e-08, 1.277078e-08, 1.498241e-07, -6.474124e-09, 2.651745e-09, 
    -9.208668e-08, 9.065332e-09, 1.473757e-08, -5.017171e-09, 1.553174e-08, 
    6.284608e-10, 8.594512e-10, -8.131451e-10, -3.130792e-09, 6.877485e-10, 
    2.582169e-08, 5.058003e-08, 3.01938e-09, 1.045976e-09, -8.93408e-10, 
    -2.697618e-09, 5.84879e-09, 3.641276e-09, 2.645922e-08, 1.571499e-08, 
    5.813945e-10, -1.231938e-08, 1.564885e-09, 9.001481e-08, 2.385661e-09, 
    -2.228381e-08, -2.227428e-08, 1.949326e-08, -1.061204e-08, -2.052445e-09, 
    -2.124011e-09, 1.810371e-09, -1.985537e-09, -5.091394e-10, 1.708202e-09, 
    -5.197762e-09, 3.784123e-09, 1.000672e-09, 7.887593e-10, 5.001084e-10, 
    -3.421405e-09, -1.712124e-10, -1.314845e-09, -2.132623e-08, 
    -7.728033e-09, 4.517005e-10, 2.723652e-10, -2.492229e-12, -2.302514e-11, 
    5.750508e-09,
  -6.282335e-09, -3.583978e-10, 2.684942e-09, 3.063462e-09, 2.597744e-11, 
    -1.828653e-10, -6.744585e-09, -8.014297e-09, -5.989477e-09, 
    -1.214357e-08, -3.804757e-09, 4.948276e-09, 5.152856e-10, 1.144883e-09, 
    3.293729e-08, -4.808874e-09, -2.728285e-08, 8.691131e-09, -3.267753e-08, 
    -4.262517e-09, 1.329465e-08, 5.824973e-09, 6.412279e-09, 6.240782e-09, 
    -5.895231e-10, -1.130559e-09, 1.483613e-11, -1.580958e-08, -2.12321e-08, 
    9.981846e-08, -3.992233e-08, -7.669939e-09, -2.578707e-08, 4.875784e-08, 
    9.56345e-09, 4.768214e-08, 5.31349e-09, 8.492833e-10, -3.009205e-08, 
    -1.250684e-08, 6.975514e-08, 3.1784e-09, 5.360732e-09, -1.194677e-08, 
    -1.710561e-08, -1.39127e-07, -5.788985e-08, 6.218596e-08, -3.054879e-09, 
    1.274714e-11, 7.323919e-10, -6.984408e-09, 2.987765e-08, -2.517481e-10, 
    9.589299e-09, -1.083151e-10, -6.770358e-08, -3.945286e-09, -9.3666e-08, 
    5.469314e-08, -1.943476e-09, -2.019306e-09, -2.097067e-09, 2.802813e-09, 
    1.022444e-08, 2.399099e-08, 4.38269e-08, 8.851089e-08, -3.282622e-08, 
    2.464219e-09, -1.230138e-07, -2.504288e-08, 1.406977e-08, -3.348248e-09, 
    1.817523e-08, 1.703256e-09, 6.469492e-10, -1.343679e-09, -3.832848e-09, 
    -7.268568e-10, 2.533724e-08, 7.686911e-08, 3.654463e-09, -1.698481e-10, 
    -3.592277e-09, 8.347456e-10, 1.899821e-09, 7.457686e-09, 6.678655e-08, 
    1.770806e-08, -3.495359e-09, -4.396583e-08, 7.013057e-11, 2.004373e-08, 
    -2.939885e-09, -2.28551e-08, -3.430156e-08, 4.656488e-08, -1.405783e-08, 
    -3.684295e-09, 1.460023e-09, 7.704628e-10, -3.232472e-09, -1.258599e-09, 
    4.567937e-10, -6.749417e-09, 4.142009e-09, 8.962388e-09, 1.33025e-09, 
    1.479066e-10, -2.483489e-09, -2.572165e-10, -2.278512e-09, -1.810832e-08, 
    5.89813e-09, 5.117897e-10, 6.284608e-10, -1.170619e-11, 6.074785e-11, 
    6.481116e-09,
  -3.254911e-09, -4.484377e-10, -3.51389e-09, 2.494284e-08, -4.714025e-10, 
    -2.999627e-10, -4.013316e-09, -1.040149e-08, 1.560562e-08, -1.387832e-09, 
    7.210986e-09, 5.423374e-09, -3.156515e-10, 1.322746e-10, 5.504432e-09, 
    -1.013053e-08, -3.33387e-08, 9.438509e-09, -3.878e-08, 3.307719e-10, 
    7.799542e-09, -1.573841e-08, -8.935956e-09, 3.923503e-09, -7.605081e-10, 
    -4.858691e-09, 9.80549e-11, -1.850896e-08, -4.606824e-08, 1.171529e-07, 
    -6.355555e-08, 1.346831e-08, -2.287544e-08, 2.996836e-08, 2.303983e-08, 
    3.650899e-08, 8.103427e-09, 1.316977e-09, -1.171486e-09, -3.236971e-08, 
    7.580417e-08, 3.488537e-09, 1.101458e-08, 3.67692e-09, 7.615483e-09, 
    -1.439468e-07, -3.871378e-08, 5.784295e-08, -2.271576e-08, 3.594991e-10, 
    3.710284e-09, -5.242833e-08, 2.897674e-08, 1.119827e-09, 1.225789e-08, 
    -3.834657e-10, -6.200202e-08, 1.453929e-08, -1.199755e-07, 5.320483e-08, 
    -2.741274e-09, -2.340187e-09, 6.412506e-10, -6.666607e-09, 1.510333e-08, 
    1.391584e-09, 4.039663e-08, 1.168456e-08, -4.227371e-08, -7.609117e-09, 
    -9.253944e-08, -2.225232e-08, 2.794934e-09, 1.82564e-09, 1.770891e-08, 
    2.858144e-09, -2.367528e-10, -6.164328e-09, -4.26376e-09, -1.054445e-10, 
    3.242963e-08, 1.121734e-07, 3.549758e-09, -2.82256e-09, -4.446861e-10, 
    6.804328e-09, 1.878442e-08, 8.099676e-09, 1.174242e-07, 4.702707e-08, 
    -6.155972e-09, -8.292274e-08, -1.509818e-09, -2.009498e-07, 
    -4.633364e-09, -6.755094e-08, -4.635286e-08, 6.881368e-08, -1.68024e-08, 
    -6.757034e-09, 2.174659e-09, -1.117613e-10, -4.715439e-09, 1.221949e-09, 
    -9.859491e-10, -1.094628e-08, 4.076298e-09, 2.245639e-08, 4.406218e-09, 
    1.572914e-09, -9.95044e-10, 6.535288e-10, -1.696492e-09, -1.021709e-08, 
    8.225186e-09, 6.118966e-10, 1.122928e-09, -6.44107e-12, 1.366516e-10, 
    7.281926e-09,
  -1.041872e-08, -4.00405e-10, -3.626269e-09, 6.633741e-08, -4.009735e-09, 
    -7.163408e-10, -3.000082e-09, -6.924552e-09, 1.77871e-08, 1.544959e-08, 
    1.404203e-08, 2.000888e-09, -1.191438e-10, 4.584876e-09, -1.70769e-09, 
    -1.072848e-08, -4.447387e-08, 1.401287e-08, -4.798365e-08, 1.237595e-08, 
    -1.038848e-08, -2.181753e-08, -2.383081e-08, -8.638153e-09, 
    -5.844413e-09, -9.328573e-09, 3.23696e-08, -1.674402e-08, -3.346895e-08, 
    6.508401e-08, -6.782113e-08, 1.345074e-08, -1.312935e-08, 6.565415e-09, 
    3.632374e-08, 1.708906e-08, 8.834661e-09, 1.733596e-09, 1.951275e-08, 
    -5.138218e-08, 9.13478e-08, 3.979039e-09, 1.540784e-08, 8.528113e-09, 
    6.677851e-09, -1.122471e-07, -6.008236e-09, 3.821168e-08, -5.915328e-08, 
    8.821246e-10, 9.824944e-09, -9.836356e-08, 1.928342e-08, 7.69062e-09, 
    1.358092e-08, -4.208687e-10, -4.769959e-08, 3.252534e-09, -9.421588e-08, 
    4.100885e-08, 5.336233e-09, -8.873258e-10, 2.464049e-09, -1.881374e-08, 
    2.310976e-08, 1.967419e-08, 3.248897e-08, 4.754725e-09, -1.275487e-08, 
    -3.712387e-08, -2.713136e-08, 6.976052e-09, -2.022591e-08, 1.597414e-09, 
    1.187675e-08, 3.803848e-09, -5.270238e-10, -1.243816e-08, -4.323818e-09, 
    -1.234639e-10, 3.242792e-08, 1.393943e-07, 2.364288e-09, -3.832952e-09, 
    1.829221e-09, 8.769121e-09, 2.448462e-08, 5.745505e-09, 1.543677e-07, 
    1.046806e-07, -6.700702e-09, -1.161716e-07, -1.443681e-09, -3.646351e-07, 
    5.233346e-09, -9.819323e-08, -5.743075e-08, 2.429877e-07, -2.025752e-08, 
    -1.001538e-08, -1.236685e-09, 2.200764e-10, -4.512891e-09, 9.419452e-10, 
    1.429726e-09, -3.486059e-08, 8.891448e-10, 2.750312e-08, 1.053149e-08, 
    2.051138e-09, 4.963567e-10, 1.240323e-09, -6.754135e-10, -1.090484e-09, 
    2.393222e-09, 7.438644e-10, 1.426429e-09, -7.386802e-11, 2.098304e-10, 
    1.066189e-08,
  -2.118304e-08, 1.455192e-11, 4.3201e-12, 9.775158e-08, -6.97105e-09, 
    -1.089802e-09, 3.119339e-09, -1.721105e-09, 8.997631e-09, 1.213289e-08, 
    1.123192e-08, -1.567741e-10, -1.863327e-10, -7.881681e-09, -1.833428e-09, 
    2.714008e-08, -6.333283e-08, 1.786236e-08, -5.426307e-08, 2.664524e-08, 
    -4.208107e-08, -1.245053e-08, -1.135265e-08, -8.353823e-09, 
    -5.054972e-09, -2.500997e-09, 1.066644e-08, -2.66665e-08, -5.363518e-09, 
    -5.35681e-09, -4.673745e-08, 1.585666e-07, -1.959256e-08, -2.437184e-08, 
    6.64885e-08, -1.741455e-08, 9.673794e-09, 1.636451e-09, 2.744719e-08, 
    -6.740925e-08, 1.186811e-07, 2.198476e-09, 1.610917e-08, 1.353858e-08, 
    -2.154638e-08, -1.039522e-07, 1.934461e-08, 8.876839e-09, -9.586272e-08, 
    -1.32701e-10, 9.95243e-10, -9.973837e-08, -1.989316e-08, 1.255007e-08, 
    1.316975e-08, -4.337153e-10, -3.081573e-08, -1.637333e-08, -3.103377e-08, 
    3.760702e-08, 8.307893e-09, -3.007017e-10, 3.67254e-09, -3.234868e-08, 
    2.755633e-08, -3.258549e-08, 2.193019e-08, 1.080321e-08, 6.542336e-09, 
    -2.794104e-08, -1.031367e-09, 1.844967e-08, -3.249727e-08, -1.040689e-09, 
    1.947978e-09, 3.820446e-09, -1.369443e-09, -1.760657e-08, -3.731304e-09, 
    1.245894e-09, 3.741809e-08, 1.846192e-07, 1.055412e-09, -1.933699e-09, 
    2.413685e-09, -1.165643e-08, 5.572247e-09, 1.293756e-09, 1.946356e-07, 
    1.783895e-07, -4.538265e-09, -1.254853e-07, -6.95195e-10, -4.342947e-07, 
    1.469357e-08, -3.450377e-07, -6.299922e-08, 1.541816e-07, -1.994692e-08, 
    -1.237822e-08, -3.694515e-08, 3.449458e-09, 8.554395e-09, 1.502507e-09, 
    2.147601e-08, -6.493269e-08, -1.712874e-08, 3.625416e-08, 1.997216e-08, 
    -1.242029e-09, -1.757485e-09, 1.126637e-09, -3.328751e-10, 2.866045e-09, 
    7.484005e-10, 9.43794e-10, 1.569688e-09, -3.669065e-10, 2.547651e-10, 
    2.03197e-08,
  -1.728313e-08, 4.351932e-10, 4.433787e-11, 8.005702e-08, -2.267097e-08, 
    2.710863e-09, 8.625648e-09, -4.256663e-09, 8.895199e-09, 1.486342e-09, 
    -1.917329e-09, -3.86774e-09, 1.804779e-09, -4.654555e-08, -5.344305e-09, 
    6.754349e-08, -8.943357e-08, 2.039371e-08, -5.193969e-08, 2.88411e-08, 
    -5.765412e-08, -8.509232e-09, -4.43174e-09, -2.163233e-09, 1.324224e-09, 
    6.349069e-09, 6.689936e-08, -2.261856e-08, 3.91185e-09, -2.560114e-09, 
    -4.134859e-08, 1.096266e-07, 9.764562e-10, -7.006781e-08, 1.048205e-07, 
    -7.219285e-08, 1.217279e-08, 1.650989e-09, 3.122261e-08, -8.599865e-08, 
    1.479377e-07, 1.569447e-09, 1.82157e-08, 1.358934e-08, -1.664432e-08, 
    -1.060323e-07, 2.87925e-08, -2.610258e-08, -1.174505e-07, -3.015479e-09, 
    1.047081e-08, -9.937321e-08, -3.602005e-08, 1.215792e-08, 9.49569e-09, 
    -8.017196e-10, -2.281843e-08, -2.780938e-08, 2.403875e-08, 3.854004e-08, 
    3.426521e-09, -2.080469e-10, 8.006623e-09, -3.947569e-08, 2.434306e-08, 
    -4.43406e-08, 8.546749e-09, 3.770833e-08, 1.422529e-08, -2.021386e-08, 
    -8.990469e-09, 3.203286e-08, -1.237208e-08, -4.412641e-09, -1.039568e-08, 
    1.559556e-09, -1.189122e-09, -1.97289e-08, -2.467343e-09, -7.809717e-09, 
    4.462686e-08, 2.057876e-07, 1.523915e-09, 1.226681e-10, -9.83232e-09, 
    -1.628803e-08, -8.82892e-09, -2.061256e-09, 2.171996e-07, 2.461458e-07, 
    -7.117933e-10, -9.692523e-08, -1.299469e-09, -4.581457e-07, 1.851345e-08, 
    -6.336585e-07, -7.122308e-08, 1.235742e-08, -1.70694e-08, -1.474127e-08, 
    -9.096084e-08, 2.359144e-09, -1.033563e-09, 1.640046e-09, 1.294063e-08, 
    -7.951292e-08, -3.385253e-08, 3.410048e-08, 3.336663e-08, -2.715069e-09, 
    -8.352572e-09, -1.458261e-09, -3.111609e-10, -1.210651e-09, 4.433673e-09, 
    9.177825e-10, 1.945324e-09, -4.682796e-10, 2.329799e-10, 3.571006e-08,
  -7.046253e-09, 2.907541e-10, 2.177103e-11, 9.824191e-09, -3.879785e-08, 
    8.083759e-09, 1.216966e-08, -5.131085e-09, 1.868159e-09, 2.162153e-09, 
    -1.87714e-09, -4.638366e-09, 3.426237e-09, -4.849829e-08, -1.400002e-08, 
    1.041135e-07, -1.264062e-07, 2.098443e-08, -4.117986e-08, 1.943812e-08, 
    -3.556733e-08, -2.056782e-08, -5.417178e-11, -3.839261e-09, 2.686704e-09, 
    2.243894e-09, -2.930454e-08, -2.45779e-08, -2.818564e-08, 1.982761e-08, 
    -4.063162e-08, 7.381499e-08, 1.248139e-08, -8.558953e-08, 9.162721e-08, 
    -1.221475e-07, 1.355862e-08, 1.511808e-09, 4.072052e-08, -1.069299e-07, 
    1.444136e-07, 5.047866e-09, 1.670247e-08, 1.341882e-08, 2.771407e-08, 
    -9.266074e-08, 2.53151e-08, -5.743681e-08, -1.252893e-07, -6.486339e-09, 
    2.451341e-08, -1.325802e-07, -2.315915e-08, 7.906113e-09, 4.201496e-09, 
    -8.916459e-10, -1.614859e-08, -3.715609e-08, 8.908827e-08, 3.69445e-08, 
    -2.35417e-09, -2.156071e-10, 1.92353e-08, -3.700758e-08, 1.367404e-08, 
    -6.7244e-08, -8.581139e-09, 5.817412e-09, -1.784821e-08, -2.111261e-08, 
    -3.83846e-08, 5.041539e-08, 7.049096e-09, -8.173345e-09, -1.064651e-08, 
    -5.082882e-09, -1.226738e-09, -2.213224e-08, -4.482644e-10, 
    -8.996778e-09, 4.905473e-08, 1.964139e-07, 4.440778e-09, -1.830927e-10, 
    -1.323491e-08, -4.206294e-08, -7.536465e-08, 2.154309e-09, 2.288849e-07, 
    2.955974e-07, 2.226159e-09, -4.982404e-08, -9.278835e-10, -3.36936e-07, 
    2.340465e-08, -8.394136e-07, -9.234369e-08, -4.23546e-09, -1.147924e-08, 
    -1.705008e-08, -9.157321e-08, -1.237938e-08, -2.376755e-08, 1.65317e-09, 
    -1.21168e-08, -6.234319e-08, -2.197766e-08, 2.816347e-08, 5.100657e-08, 
    1.358387e-09, -8.263726e-09, -4.21943e-09, 5.196057e-10, -5.51421e-09, 
    6.153925e-09, 2.776574e-10, 2.330452e-09, -5.149658e-10, 1.815508e-10, 
    4.332168e-08,
  3.596313e-09, 3.144009e-10, -9.147868e-09, -4.489522e-08, -2.286964e-08, 
    1.940674e-08, 1.442612e-08, 1.498222e-09, -6.228277e-09, -9.843745e-09, 
    -3.689649e-09, -1.408182e-09, 2.177615e-09, 3.783441e-09, -2.616201e-08, 
    1.263407e-07, -1.596917e-07, 2.052298e-08, -6.182262e-09, -2.11358e-08, 
    2.805166e-09, -3.77284e-08, 6.722871e-10, -1.048818e-09, 1.937394e-09, 
    -5.671097e-09, -2.790131e-08, 3.291234e-11, -2.520227e-08, 3.066071e-08, 
    -3.021427e-08, 8.747855e-08, -5.492723e-09, 3.640309e-09, 1.025484e-08, 
    -1.63003e-07, 1.463253e-08, 7.764527e-10, 5.970668e-08, -1.348676e-07, 
    7.371053e-08, 7.023857e-09, 1.474547e-09, 1.442124e-08, 3.043937e-08, 
    -6.297756e-08, 1.026569e-08, -7.421198e-08, -1.05504e-07, -8.468639e-09, 
    3.217396e-08, -1.337207e-07, -3.447838e-09, 4.360811e-09, 2.352408e-10, 
    -3.453238e-10, -1.781615e-08, -4.251429e-08, 1.101907e-07, 5.933092e-08, 
    -1.491173e-09, -1.532328e-09, 2.160533e-08, -3.416507e-08, -2.556419e-09, 
    -7.791726e-08, -2.282781e-08, 2.497353e-08, -6.185365e-08, -2.845621e-08, 
    -9.908678e-08, 4.418115e-08, 4.867405e-08, 2.1451e-09, 1.833439e-09, 
    -8.271115e-09, -1.675602e-09, -2.378169e-08, 1.776954e-10, 2.573358e-09, 
    5.045166e-08, 1.942361e-07, 9.26741e-09, 1.431033e-09, 2.655156e-10, 
    -4.267707e-08, 1.121725e-07, 7.627989e-09, 2.347377e-07, 3.214166e-07, 
    -4.856133e-10, -2.193193e-08, 9.439987e-10, -2.007193e-07, 2.225778e-08, 
    -9.74131e-07, -1.354805e-07, -9.652183e-09, -6.836842e-09, -1.64482e-08, 
    4.914114e-10, -3.19024e-08, -3.272197e-08, 7.002114e-10, -8.275663e-09, 
    -4.011423e-08, -5.37824e-09, 7.769927e-10, 7.611965e-08, 1.465907e-08, 
    -2.056311e-09, -2.75935e-09, -5.088054e-10, -6.196672e-09, 3.556067e-09, 
    -6.300979e-10, 2.360579e-09, -9.043895e-10, 1.453273e-10, 3.969939e-08,
  5.192703e-09, 3.29635e-10, -5.775917e-09, -5.167107e-08, -1.530174e-08, 
    2.72849e-08, 1.773464e-08, 1.48213e-08, -1.211276e-09, -2.246509e-09, 
    -9.075052e-10, -4.508252e-10, 9.097278e-09, 5.843788e-09, -1.708219e-08, 
    1.261221e-07, -1.669618e-07, 6.906055e-08, 3.345878e-08, -9.019624e-08, 
    3.443444e-08, -4.680186e-08, 1.487081e-09, -2.943921e-10, -2.189779e-09, 
    -5.175991e-09, -2.791495e-08, 2.083306e-08, -1.992549e-08, 1.586528e-08, 
    -3.686858e-08, 5.562907e-08, -4.621995e-09, 3.314523e-08, -4.272732e-08, 
    -1.633366e-07, 1.539364e-08, 5.359482e-10, 8.688409e-08, -1.703716e-07, 
    -6.368638e-08, 7.806136e-09, -6.503086e-08, 1.256465e-08, 7.489859e-09, 
    -2.805047e-08, 3.23729e-09, -6.723647e-08, -8.092642e-08, -1.016033e-08, 
    3.475451e-08, -1.030219e-07, 1.647447e-08, 8.084418e-09, -3.427658e-09, 
    -2.760885e-10, -2.761959e-08, -5.683422e-08, 8.946897e-08, 1.223404e-07, 
    2.983313e-09, -2.744457e-09, 1.579639e-08, 2.06918e-09, -2.742362e-08, 
    -5.881196e-08, -2.268388e-08, 3.822055e-08, -9.144816e-08, -3.596136e-08, 
    -1.696629e-07, 8.435961e-09, 1.515311e-07, 1.293472e-09, 8.86539e-09, 
    5.513982e-09, -2.838718e-09, -2.460439e-08, -7.589392e-10, -3.803223e-09, 
    4.632716e-08, 2.135217e-07, 1.496147e-08, 4.509218e-09, 5.449181e-09, 
    -1.774498e-08, 1.469368e-07, 1.03858e-08, 2.409459e-07, 3.301241e-07, 
    -8.776453e-09, -1.382854e-08, 1.644082e-09, -9.894923e-08, 2.575945e-08, 
    -9.822845e-07, -1.685523e-07, 1.616144e-08, -2.752984e-09, -1.216284e-08, 
    1.117167e-07, -3.084923e-08, -3.440702e-08, 9.738343e-10, 1.166467e-08, 
    -2.721998e-08, -9.66628e-09, -1.490258e-08, 8.89608e-08, 2.961775e-08, 
    8.298571e-10, 1.788123e-09, 9.933387e-10, -4.583569e-09, 9.498535e-11, 
    -1.691797e-09, 3.895252e-09, -1.392824e-09, 1.678515e-10, 2.386165e-07,
  2.387196e-09, -1.29603e-11, 2.777483e-09, -2.064644e-08, 7.590074e-09, 
    3.260061e-08, 2.378499e-08, 5.627066e-08, 1.730177e-08, -1.576109e-08, 
    1.9254e-09, -1.47395e-09, 3.91401e-09, -1.711783e-08, 2.680974e-08, 
    1.109771e-07, -1.716236e-07, 6.602903e-08, 7.381016e-08, -1.188541e-07, 
    3.834793e-08, -4.639492e-08, 6.666596e-10, 5.700258e-10, -1.584408e-08, 
    3.824539e-09, -3.169362e-09, 1.766261e-08, -2.107902e-08, -2.655156e-09, 
    -6.022606e-08, 3.952118e-08, 8.611437e-09, 3.183266e-08, -3.131117e-08, 
    -1.468472e-07, 1.376683e-08, 5.2448e-10, 1.025951e-07, -2.102082e-07, 
    -1.765655e-07, 7.926815e-09, -2.055158e-07, 2.140574e-08, -7.447625e-10, 
    -1.172077e-08, 2.756468e-08, -3.470402e-08, -6.620903e-08, -1.112714e-08, 
    3.518151e-08, -7.955271e-08, 3.214794e-08, 1.251524e-08, -7.609069e-09, 
    -1.53193e-10, -3.906473e-08, -8.211532e-08, 6.577028e-08, 2.178484e-07, 
    2.949719e-09, 7.288463e-09, 6.119421e-09, 1.997905e-08, -5.69275e-08, 
    -2.170805e-08, -2.045101e-08, 2.194247e-08, -9.899156e-08, -3.759999e-08, 
    -1.322464e-07, -4.279491e-08, 2.237115e-07, -9.448854e-09, 5.383049e-09, 
    1.353874e-08, -3.350294e-09, -2.362765e-08, -1.028224e-09, -8.356892e-09, 
    3.835186e-08, 2.369214e-07, 1.69191e-08, 1.024932e-08, -4.281446e-09, 
    2.672823e-08, 7.48098e-08, 7.493441e-09, 2.44851e-07, 3.195493e-07, 
    1.105036e-10, -1.688445e-08, 3.001617e-10, -1.34643e-08, 5.219056e-08, 
    -8.034477e-07, -1.116707e-07, 1.709498e-08, 6.734467e-09, -6.802634e-09, 
    -1.616047e-08, -9.528527e-09, -2.38113e-08, 2.427889e-09, 1.142553e-09, 
    -6.623736e-09, -5.938318e-09, -4.538606e-09, 8.174504e-08, 3.072216e-08, 
    -1.956892e-09, 5.231527e-09, 1.764079e-09, 4.868525e-09, -6.691266e-09, 
    -2.942829e-09, 3.247848e-09, -1.310028e-09, 2.008349e-10, 7.640324e-09,
  6.938876e-10, -1.967749e-09, 9.71221e-09, 1.428879e-08, 3.01672e-08, 
    2.831479e-08, 3.214899e-08, 8.402066e-08, 4.54001e-08, -7.61043e-08, 
    -1.504696e-08, -5.759205e-09, -1.138579e-08, -4.250734e-08, 4.979159e-08, 
    8.750946e-08, -1.806628e-07, 4.160762e-08, 1.970285e-07, -1.208351e-07, 
    1.43836e-08, -2.716666e-08, 2.404477e-11, 4.769163e-11, 1.110436e-09, 
    4.673001e-08, 8.903669e-09, 1.257575e-08, -2.638927e-08, -4.612104e-09, 
    -8.915941e-08, 8.732576e-08, 9.057146e-09, 4.790917e-08, -1.892317e-10, 
    -1.452661e-07, 1.095976e-08, -1.289294e-09, 1.004154e-07, -2.457916e-07, 
    -2.030532e-07, 6.001244e-09, -2.761565e-07, 3.13494e-08, -1.007635e-08, 
    2.282553e-08, 4.411334e-09, -9.877112e-09, -5.587236e-08, -1.747708e-09, 
    3.207174e-08, -7.683644e-08, 4.014347e-08, 1.88304e-08, -1.263605e-08, 
    2.563638e-11, -5.989529e-08, -9.930874e-08, 3.764468e-08, 3.083519e-07, 
    -1.330648e-09, -1.109385e-08, -1.988434e-08, 5.605523e-09, -8.016264e-08, 
    -2.261396e-08, -1.757331e-08, -1.87157e-09, -9.416368e-08, -2.678627e-08, 
    -1.260474e-08, -6.854071e-08, 9.745071e-08, -6.722587e-09, 9.01681e-09, 
    4.770698e-09, 4.036167e-10, -1.548131e-08, -1.062187e-09, -2.292842e-08, 
    3.047938e-08, 2.415411e-07, 1.537836e-08, 2.54542e-08, -1.317545e-08, 
    9.281365e-08, 4.088332e-08, 2.942613e-09, 2.483391e-07, 2.906324e-07, 
    8.32955e-09, -2.894159e-08, -1.822457e-09, 6.164095e-08, 8.435376e-08, 
    -5.081941e-07, -1.325839e-07, -3.670567e-08, 1.35953e-08, -1.799174e-09, 
    -3.5364e-09, 8.310792e-09, -1.835843e-08, 3.394845e-09, -4.068926e-08, 
    -5.720591e-08, 1.033129e-09, 1.46087e-08, 5.884243e-08, 1.816915e-08, 
    -4.754895e-09, 3.414641e-09, 2.121112e-09, 1.285042e-08, -1.332825e-08, 
    -3.311868e-09, 3.33435e-09, -1.094392e-09, 2.322906e-10, -5.093858e-08,
  1.473211e-09, -8.003838e-09, 1.090183e-08, 4.713974e-08, 7.341026e-08, 
    3.182203e-08, 2.724533e-08, 6.029205e-08, 5.406156e-08, -5.987812e-08, 
    -6.309023e-08, 8.929095e-08, -1.214977e-08, -3.644737e-08, 1.965412e-08, 
    7.024695e-08, -1.97684e-07, -1.543071e-09, 3.949292e-08, -1.321991e-07, 
    1.112028e-09, 1.104326e-08, -4.999322e-09, -1.634004e-08, 7.698247e-09, 
    2.576661e-08, 2.824606e-09, 5.786831e-09, -3.536474e-08, -3.842916e-08, 
    -8.513365e-08, 7.908005e-08, -1.468777e-09, 2.395001e-08, 2.330631e-08, 
    -1.726067e-07, 9.589496e-09, -1.277087e-09, 8.621754e-08, -2.761543e-07, 
    -1.822472e-07, 1.254818e-09, -2.11991e-07, 2.605586e-08, -2.143105e-08, 
    4.126053e-08, -1.804608e-09, -7.479883e-09, -4.949221e-08, 7.792991e-09, 
    2.448867e-08, -8.633145e-08, 4.517545e-08, 1.903955e-08, -1.710671e-08, 
    -2.830802e-11, -9.412128e-08, -1.176162e-07, 2.411529e-08, 3.485969e-07, 
    -4.268315e-09, -2.357592e-07, 8.0549e-08, 4.666855e-08, -1.04989e-07, 
    -2.674136e-08, -1.154712e-08, -1.840471e-08, -8.092576e-08, 
    -1.779341e-08, 4.359691e-08, -3.810948e-08, 2.459973e-08, -4.009678e-09, 
    1.72148e-08, -6.945697e-10, 5.531007e-09, -1.190344e-08, -2.949378e-09, 
    -5.481769e-08, 2.239545e-08, 2.340236e-07, 1.000939e-08, -3.680117e-08, 
    -3.942586e-08, 8.556725e-08, -1.37855e-07, 6.564846e-10, 2.470113e-07, 
    2.634343e-07, 1.139091e-08, -4.235968e-08, -2.965351e-09, 1.069951e-07, 
    7.883654e-08, -3.606723e-07, -1.559519e-07, -6.0368e-08, 2.114786e-08, 
    -1.954606e-09, 3.4675e-08, 1.05943e-08, -1.935368e-08, 7.946788e-09, 
    2.834832e-08, -6.957822e-08, 2.362356e-09, 1.610732e-08, 2.729331e-08, 
    1.509932e-09, -1.420921e-08, -4.83567e-10, -1.305693e-10, 1.075051e-08, 
    -9.307257e-09, -2.918034e-09, 3.389928e-09, -1.100585e-09, 3.174065e-10, 
    -9.232411e-08,
  2.732236e-09, -1.549768e-08, 3.486775e-10, 3.300954e-08, 6.029643e-08, 
    3.468301e-08, 1.9916e-08, 4.413448e-08, 6.358994e-08, -3.266985e-08, 
    -6.370453e-08, 3.911554e-07, -1.198225e-08, -2.137028e-08, -3.542038e-08, 
    5.469044e-08, -2.22626e-07, -1.222668e-08, -1.380107e-08, -8.604172e-08, 
    -9.061398e-08, 3.750387e-07, 1.431789e-07, -3.516164e-07, 4.65908e-08, 
    1.260025e-08, -2.807042e-09, 5.076458e-09, -6.754419e-08, -6.36486e-08, 
    -3.601679e-08, 3.630487e-08, -2.071295e-08, 6.840639e-08, 2.505942e-08, 
    -2.202847e-07, 1.07387e-08, -1.303334e-09, 6.751532e-08, -3.011087e-07, 
    -1.251146e-07, -1.623108e-07, -4.873385e-08, 3.575984e-08, -3.515709e-08, 
    1.206706e-08, -6.386108e-08, -3.068914e-08, -5.524755e-08, 1.618022e-08, 
    2.873861e-09, 7.993856e-08, 5.31297e-08, 1.626524e-08, -2.07499e-08, 
    -1.180069e-10, -8.48728e-08, -1.338116e-07, 2.470651e-08, 3.424262e-07, 
    -2.361617e-09, -3.76732e-08, -4.076799e-08, 6.167509e-08, -1.194639e-07, 
    -2.576814e-08, 1.058049e-08, -3.256343e-08, -6.155335e-08, -3.679247e-09, 
    8.453151e-08, 2.935678e-08, 4.527385e-08, -1.062961e-08, -1.623021e-08, 
    -6.237428e-09, 4.896208e-10, -4.726303e-09, -6.110986e-09, -6.151174e-08, 
    6.304958e-09, 2.271329e-07, 2.911293e-09, -2.07807e-08, -6.422931e-08, 
    2.184981e-08, -1.175848e-07, -9.476366e-09, 2.30583e-07, 2.465871e-07, 
    1.910246e-08, -5.110831e-08, -7.053018e-09, 1.234571e-07, 8.049835e-08, 
    -2.765692e-07, -1.326081e-07, -7.170536e-08, 3.099115e-08, 4.342339e-08, 
    1.070426e-07, 6.154011e-10, -2.309845e-08, 1.589369e-08, -4.891615e-08, 
    -7.854635e-08, -1.640581e-08, 3.113314e-09, -7.268113e-09, -2.123386e-08, 
    -2.924855e-08, 1.905505e-09, -5.708216e-10, 1.476189e-08, -3.698119e-09, 
    -1.494823e-09, 5.41641e-09, -9.945609e-10, 4.077236e-10, -6.451444e-08,
  2.76026e-09, -2.017606e-08, -2.96605e-08, -2.819036e-09, 6.948937e-09, 
    1.559255e-08, 1.793427e-08, 4.246425e-08, 7.609805e-08, -1.588529e-08, 
    2.821679e-08, 2.199126e-07, 1.233474e-08, -1.852487e-08, -6.856914e-08, 
    6.420977e-08, -2.453727e-07, 2.197947e-08, 2.699664e-09, -7.743625e-08, 
    -1.150811e-07, -3.917017e-08, -9.704928e-08, 6.43783e-08, 8.316027e-08, 
    -7.161867e-08, 4.602896e-09, 1.089751e-08, -4.556188e-08, -6.953707e-08, 
    -4.503505e-08, -1.718428e-08, -5.460112e-08, 5.159831e-08, 1.269581e-08, 
    -2.717027e-07, 1.869865e-08, -1.645844e-09, 4.906923e-08, -2.99673e-07, 
    -5.699017e-08, -4.136319e-08, 2.092008e-09, 3.314526e-08, -3.264478e-08, 
    -4.874488e-08, -8.407102e-08, -6.268289e-08, -1.74589e-08, 1.951972e-08, 
    5.082427e-09, -1.059944e-07, 6.057102e-08, 2.004766e-08, -2.303872e-08, 
    -3.449827e-10, -1.096907e-09, -1.467107e-07, 3.2734e-08, 3.536606e-07, 
    -3.961418e-10, 2.529413e-08, -7.006958e-08, 9.523168e-08, -1.206829e-07, 
    -2.082157e-08, 1.510002e-07, -3.75606e-08, -3.591441e-08, 1.89379e-08, 
    1.022262e-07, 7.534408e-08, 4.062912e-08, -3.024053e-08, -1.499579e-08, 
    -7.954498e-09, -7.397659e-09, 4.527408e-09, -9.359451e-09, -1.691143e-08, 
    -1.039376e-08, 2.142393e-07, -2.164029e-10, 6.602198e-08, -5.139924e-08, 
    1.257055e-07, -1.154093e-07, -1.744803e-08, 1.977866e-07, 2.26141e-07, 
    -1.691484e-08, -4.994937e-08, -3.763375e-09, 1.074735e-07, 6.929798e-08, 
    -2.867854e-07, -1.172349e-07, 4.417956e-08, 3.47531e-08, 1.32451e-07, 
    2.743206e-07, -1.765942e-08, -2.659927e-08, 2.487454e-08, -7.487989e-08, 
    -5.595172e-08, -3.565788e-10, -7.976098e-09, -3.213205e-08, 
    -4.028203e-08, -3.040583e-08, 1.023335e-08, 4.39735e-09, 2.560813e-08, 
    -2.590525e-09, -2.208367e-10, 6.520821e-09, -8.602612e-10, 4.925766e-10, 
    -3.471206e-08,
  -2.831939e-10, -1.503383e-08, -6.763764e-08, -6.155631e-08, -4.459218e-08, 
    3.807941e-09, 5.208005e-08, 5.823597e-08, 7.030201e-08, 1.465537e-09, 
    7.025903e-08, -2.907143e-08, 3.389584e-08, -1.674823e-08, 3.470552e-08, 
    7.679694e-08, -2.661473e-07, 8.889742e-09, 5.967877e-08, -8.102813e-08, 
    -2.123841e-08, -1.825845e-08, -7.198912e-08, 9.623352e-08, -1.587599e-07, 
    -2.084081e-07, -4.56547e-08, 1.542901e-08, -1.291926e-08, -7.283654e-08, 
    -5.470008e-08, -4.070841e-08, -3.474213e-08, -2.537388e-08, 1.892715e-08, 
    -3.009756e-07, 1.916926e-08, -1.209884e-09, 2.89491e-08, -2.552001e-07, 
    -1.241906e-07, 1.847467e-07, -5.30153e-08, 2.480992e-08, -2.002855e-08, 
    -7.985625e-08, -7.645167e-08, -8.997472e-08, -3.224752e-08, 1.736247e-08, 
    1.392436e-09, -1.929226e-07, 7.811989e-08, 2.848321e-08, -2.628254e-08, 
    -2.409706e-09, 4.976766e-08, -1.523392e-07, 5.372835e-08, 3.831174e-07, 
    2.100592e-09, 9.832308e-08, 1.079751e-07, 9.359176e-08, -1.109937e-07, 
    -1.68726e-08, 8.184327e-08, -3.776211e-08, -1.899241e-08, 3.070443e-08, 
    1.080422e-07, 8.724021e-08, 2.385036e-09, -4.482615e-08, -1.210572e-08, 
    -8.389975e-09, 7.332687e-09, 1.723606e-09, 9.690864e-09, 1.447091e-07, 
    -2.509216e-08, 1.917626e-07, 1.046055e-08, 1.72122e-07, -1.453725e-08, 
    -4.123763e-09, -1.602722e-07, -1.189289e-08, 1.629141e-07, 1.908235e-07, 
    -1.062421e-07, -4.413052e-08, -9.908035e-09, 7.693117e-08, 1.135658e-07, 
    -3.44646e-07, -5.284858e-08, 1.04443e-08, 3.146204e-08, 5.044133e-08, 
    5.971026e-08, -4.352295e-08, -3.060637e-08, 2.596261e-08, -4.312028e-09, 
    5.283368e-09, -3.705168e-09, -2.003719e-08, -4.791207e-08, -4.860533e-08, 
    -2.561649e-08, 1.775118e-08, 1.103592e-08, 4.599121e-08, 6.678306e-09, 
    9.047653e-10, 6.299189e-09, -9.720367e-10, 5.134666e-10, -3.270145e-08,
  2.847457e-09, 7.996107e-09, -7.202124e-08, -7.471107e-08, -4.556995e-08, 
    -2.283758e-08, 1.532881e-07, 8.730427e-08, 4.698751e-08, 7.250907e-08, 
    3.836323e-08, -1.243358e-07, 5.957742e-08, 1.033612e-07, -1.060818e-07, 
    8.774858e-08, -2.645752e-07, -2.38623e-09, 1.378319e-08, -1.495889e-07, 
    6.131933e-08, 1.602581e-08, -3.221515e-08, 2.046869e-08, -1.025014e-07, 
    -2.36261e-07, -7.382772e-08, 1.568861e-08, -5.165873e-09, -7.332864e-08, 
    -7.459329e-08, -6.139584e-08, -8.115819e-09, -4.258339e-08, 3.664542e-08, 
    -2.264516e-07, 6.962898e-09, -1.077723e-09, 1.040081e-08, -1.917614e-07, 
    -1.098923e-07, 1.967947e-07, -9.097147e-08, 1.499126e-08, -2.589189e-08, 
    -7.967668e-08, -8.071248e-08, -1.641956e-07, -3.273038e-08, 1.141264e-08, 
    2.912515e-09, -1.118719e-07, 9.598426e-08, 3.451402e-08, -3.342128e-08, 
    -1.200425e-08, 6.905981e-08, -1.558466e-07, 2.173777e-07, 3.70702e-07, 
    5.912909e-09, -1.964679e-09, -1.061647e-08, 5.210269e-08, -8.204169e-08, 
    -1.42922e-08, -4.324301e-08, -4.036787e-08, -2.080282e-08, 2.406188e-08, 
    9.58949e-08, 6.404144e-08, -6.512727e-08, -4.085604e-08, -3.321736e-09, 
    -6.359812e-09, 1.000927e-09, -2.808349e-09, 2.30736e-08, 2.066666e-07, 
    -2.429641e-08, 1.685738e-07, -3.348703e-09, -3.00326e-08, 1.908012e-08, 
    -3.179315e-08, -1.595167e-07, -7.173071e-10, 1.499082e-07, 1.499166e-07, 
    -2.452788e-08, -3.537519e-08, -9.690837e-09, 4.636964e-08, 2.102684e-07, 
    -4.061815e-07, 3.208021e-08, 1.083964e-08, 2.877738e-08, -2.886672e-08, 
    -5.600839e-09, 5.434448e-08, -3.339829e-08, 2.036067e-08, 4.38402e-08, 
    3.168185e-08, 4.034803e-09, -3.066106e-08, -6.195017e-08, -5.084934e-08, 
    -2.477731e-08, 1.831341e-08, -5.006029e-09, 5.020757e-08, -2.111108e-09, 
    1.522505e-09, 8.212282e-09, -2.084718e-09, -6.609753e-10, -4.173097e-08,
  1.73722e-08, 4.309726e-08, -3.51834e-08, -3.599035e-08, -7.140972e-08, 
    -2.135009e-07, 1.159729e-07, 9.639217e-08, 4.546945e-08, -1.018012e-07, 
    -3.116435e-08, -1.037626e-07, 1.012001e-07, -1.092622e-07, -1.465998e-07, 
    9.165424e-08, -2.163698e-07, -4.379621e-08, -2.064922e-09, -6.297768e-08, 
    2.757866e-08, 1.334382e-08, 4.250074e-08, -8.176528e-09, 2.966459e-08, 
    -1.326031e-07, -2.193184e-08, 1.595055e-08, 7.234291e-09, -6.668319e-08, 
    -4.256498e-08, -4.428563e-08, -1.935581e-08, -2.790483e-08, 1.93482e-07, 
    -1.94562e-07, -1.277453e-09, -8.033822e-10, -4.162132e-09, -1.183612e-07, 
    -1.262909e-07, 1.529463e-07, -1.075975e-07, -2.266507e-10, -2.881296e-08, 
    -8.150545e-08, -7.608025e-08, -2.10405e-07, -2.527378e-08, 5.700734e-09, 
    -1.579721e-09, -8.74283e-08, 1.188276e-07, 4.171287e-08, -4.502795e-08, 
    2.46132e-11, 6.267391e-08, -1.800304e-07, 3.209283e-07, 2.394107e-07, 
    9.063859e-08, -1.176608e-08, 8.517492e-08, 4.083214e-08, -3.238331e-08, 
    -7.567735e-09, -1.243336e-07, -4.334009e-08, -2.380483e-08, 8.814652e-09, 
    7.345926e-08, 7.038523e-09, -1.218124e-07, -1.564575e-08, 9.890293e-10, 
    -7.12663e-09, -1.310309e-08, 1.195258e-08, 2.191436e-09, 2.422547e-08, 
    -1.635459e-08, 1.316511e-07, -1.174783e-08, -2.712551e-08, 4.175541e-08, 
    8.565127e-08, -1.351942e-07, 6.720597e-10, 1.36215e-07, 1.106754e-07, 
    8.751653e-08, -2.553137e-08, -1.053115e-08, 3.689988e-08, 2.738917e-07, 
    -4.557425e-07, 4.086659e-08, -2.872292e-08, 7.380947e-09, -9.100464e-08, 
    4.433497e-08, -4.705824e-08, -3.426107e-08, 1.401646e-08, 1.119842e-07, 
    3.869337e-08, 1.518339e-08, -3.936367e-08, -7.169814e-08, -5.153919e-08, 
    -2.697465e-08, -3.888658e-10, -1.924485e-08, 1.736424e-08, 9.998189e-10, 
    2.62803e-09, 7.535562e-09, -2.033325e-09, -5.27919e-10, -3.842746e-08,
  3.271549e-08, 6.997544e-08, 7.222013e-09, -1.711243e-08, -4.825117e-07, 
    -3.054226e-07, 1.102495e-08, -8.284303e-09, 7.08468e-09, -5.20443e-08, 
    -6.638624e-08, -5.958651e-08, -7.365787e-08, -9.850493e-08, 
    -1.781047e-07, 8.684076e-08, -1.642146e-07, 2.878323e-09, -7.672199e-09, 
    -3.29963e-08, -7.963564e-08, -6.91665e-09, 1.903248e-07, 6.455792e-08, 
    1.110744e-07, -5.862199e-08, -4.095358e-08, 1.606628e-08, -2.082004e-09, 
    -5.078431e-08, -3.452868e-08, -2.497057e-08, -1.340487e-08, 
    -7.066944e-09, 2.187526e-07, -2.576409e-07, -3.921127e-09, -2.434035e-10, 
    -1.465793e-08, -1.162857e-07, -1.152432e-07, 2.335343e-07, -6.136241e-08, 
    -1.731002e-08, -4.074803e-08, -7.723219e-08, -7.474426e-08, 
    -1.932022e-07, -2.847067e-08, 3.139178e-09, -1.079172e-09, 2.996973e-08, 
    1.391583e-07, 4.600335e-08, -3.611058e-08, -1.050353e-09, 5.388091e-08, 
    -1.542879e-07, 1.362179e-07, 1.407582e-07, 9.093429e-08, -7.719422e-08, 
    1.031555e-08, 3.19341e-08, 8.643809e-09, -1.296655e-09, -9.765409e-08, 
    -4.66311e-08, -1.807149e-08, -1.1201e-09, 3.583472e-08, -2.766041e-08, 
    -1.697029e-07, -1.070369e-07, 2.578646e-08, -5.194522e-09, -1.092647e-08, 
    6.091057e-09, -2.035617e-08, 1.763095e-08, -1.979362e-08, 1.27449e-07, 
    1.816886e-08, -8.843409e-08, 7.487898e-08, 8.458989e-08, -4.845293e-08, 
    -5.697814e-09, 1.406436e-07, 8.317801e-08, 7.278385e-08, -2.535177e-08, 
    -8.445653e-09, 5.798724e-08, 1.873821e-07, -4.901702e-07, 1.349814e-08, 
    -8.826504e-08, 1.528775e-08, -8.551297e-08, -1.816073e-08, 1.291296e-08, 
    -3.50952e-08, 9.212322e-09, 1.464944e-07, 2.691826e-08, 2.833491e-08, 
    -4.609598e-08, -7.991235e-08, -5.349699e-08, -2.666656e-08, 
    -5.924278e-09, -1.184861e-08, 9.185271e-09, 7.057508e-09, 4.095148e-09, 
    3.846864e-09, -1.862887e-09, -4.001777e-10, -6.750025e-08,
  3.779093e-08, 4.056341e-08, 1.137943e-08, -3.226219e-07, -5.134432e-07, 
    -1.082475e-08, 7.067399e-09, -1.612483e-08, -2.015389e-08, -2.141832e-08, 
    -7.441616e-08, -7.858677e-08, -6.1614e-08, -9.599017e-08, -1.602663e-07, 
    8.27416e-08, -7.780633e-08, 3.463657e-08, 1.520176e-08, -3.624046e-08, 
    -1.243717e-08, 4.639304e-08, 1.444465e-08, 7.708235e-08, -3.372958e-08, 
    7.719962e-09, -3.223437e-08, 7.320239e-09, -1.084055e-08, -3.487349e-08, 
    1.45464e-08, -2.577775e-08, -4.212865e-08, -1.553957e-08, 1.93989e-07, 
    -2.474559e-07, 6.34145e-11, -2.843024e-10, -2.125984e-08, -1.143778e-07, 
    -8.156755e-08, -1.443622e-07, -2.781911e-08, 1.461901e-09, -2.969267e-08, 
    -8.528269e-08, -6.105756e-08, -1.47203e-07, -1.583102e-08, 3.274145e-09, 
    2.966232e-10, -1.127694e-07, 1.505346e-07, 3.967983e-08, -2.482672e-08, 
    -1.271303e-09, 1.41083e-07, -1.324614e-07, 1.132332e-08, 1.018253e-07, 
    -4.772176e-09, -9.840511e-08, -1.406297e-07, 2.149214e-08, 4.521913e-08, 
    -4.116885e-09, -7.667956e-08, -4.321424e-08, -3.389181e-08, 
    -1.133657e-08, 3.86359e-09, -6.871613e-08, -1.751768e-07, -3.17329e-08, 
    1.854765e-09, -1.033897e-08, -8.399979e-09, 1.345711e-08, -4.472172e-08, 
    7.905982e-08, -4.586013e-08, 1.341745e-07, 3.587638e-08, -3.446718e-08, 
    8.211538e-08, -1.267478e-08, 6.340991e-08, -1.65283e-08, 1.567226e-07, 
    6.317583e-08, 8.456021e-08, -3.082822e-08, -1.976844e-09, 6.504519e-08, 
    1.198206e-07, -5.327799e-07, -1.668833e-08, -9.886236e-08, 2.496159e-08, 
    -5.330706e-08, -2.854296e-08, 5.138453e-08, -2.295887e-08, 4.79703e-09, 
    7.448915e-08, -4.526612e-09, 4.312921e-08, -5.195892e-08, -8.512922e-08, 
    -5.566488e-08, -2.706582e-08, -8.680615e-09, -3.13031e-09, 5.113236e-09, 
    7.792039e-09, 5.218078e-09, 4.293398e-09, -1.965365e-09, -2.513403e-10, 
    -1.057064e-07,
  -1.807098e-08, 1.290141e-08, -2.823695e-07, -5.550058e-07, -9.362566e-08, 
    6.369373e-08, 3.374453e-09, 1.277499e-09, -1.487786e-08, -3.950515e-08, 
    -1.055207e-07, -7.274878e-08, -8.224197e-08, 1.976002e-08, -7.061169e-08, 
    8.217289e-08, -1.857945e-08, 4.082301e-08, 4.365769e-08, -3.035564e-08, 
    3.177547e-08, -8.833354e-09, 1.772639e-08, -5.418201e-09, 2.722049e-08, 
    5.972163e-08, -5.50865e-08, 1.122908e-08, -8.870757e-08, -3.191053e-08, 
    3.394928e-08, -1.044771e-08, -4.392678e-08, -5.221352e-08, 2.854297e-07, 
    -1.732319e-07, 8.782138e-09, -7.926815e-10, -3.375828e-08, -6.874765e-08, 
    3.078728e-08, -2.641507e-07, 2.918208e-08, 7.423232e-09, -3.240757e-08, 
    -1.09689e-07, -5.598827e-08, -9.950551e-08, -2.6971e-08, 2.950948e-09, 
    1.203048e-09, -4.48656e-08, 1.451101e-07, 3.743396e-08, -2.457418e-08, 
    -1.583601e-09, 1.408221e-07, -1.414804e-07, -3.559612e-08, 1.197937e-07, 
    -1.012984e-08, 1.121138e-07, -9.937253e-08, -1.552512e-08, 5.416349e-08, 
    -7.232529e-09, -3.974799e-08, -3.306627e-08, -7.60823e-08, -2.988884e-08, 
    8.801635e-10, -9.875203e-08, -6.276821e-08, 1.094011e-07, -6.336137e-09, 
    -2.026832e-08, -1.808722e-08, 1.839044e-08, -5.463837e-08, 9.480584e-08, 
    -6.28682e-08, 1.401692e-07, 2.264812e-08, -9.081987e-09, 3.828802e-08, 
    -3.424839e-08, 1.235555e-07, -3.79099e-08, 1.147075e-07, 5.840388e-08, 
    9.097721e-08, -2.220011e-08, 6.768801e-09, 6.237245e-08, -2.488639e-08, 
    -5.940911e-07, -2.286549e-08, -7.72053e-08, 3.604589e-08, -4.543947e-08, 
    4.38414e-08, 3.499025e-09, -3.50161e-08, 4.021928e-09, 3.356524e-08, 
    -1.818989e-11, 4.963977e-08, -5.781442e-08, -8.990935e-08, -5.738684e-08, 
    -2.741967e-08, -9.517066e-09, -2.589559e-09, 4.937419e-09, 6.791197e-09, 
    6.045525e-09, 4.737998e-09, -2.002331e-09, -1.937366e-10, -8.099005e-08,
  8.556481e-08, 2.998688e-07, -2.976013e-07, -1.734023e-07, -3.717764e-08, 
    2.840011e-09, -1.333194e-08, -5.572838e-08, 1.671094e-08, -4.66672e-08, 
    -7.046788e-08, -6.965831e-08, 2.037473e-08, 4.279286e-08, 2.513434e-08, 
    8.652906e-08, -1.436898e-08, 4.574099e-08, -2.434518e-09, -4.726405e-08, 
    -1.40268e-08, -5.080324e-09, 3.980335e-08, -9.357791e-09, 1.544595e-08, 
    2.377544e-08, -7.27382e-08, 9.381552e-09, -1.293772e-07, -3.298385e-08, 
    3.098557e-08, -3.134767e-08, -2.936451e-08, -1.822661e-08, 1.054073e-07, 
    -4.792173e-08, 1.335691e-08, -8.459438e-10, -3.273374e-08, -5.516616e-08, 
    8.054458e-08, -5.100924e-08, 1.56061e-08, -1.097996e-08, -5.68408e-08, 
    -1.38314e-07, -5.2046e-08, -8.854363e-08, -3.870732e-08, 3.166654e-09, 
    2.630756e-09, -4.658841e-08, 1.286988e-07, 3.379155e-08, -2.216644e-08, 
    -4.736421e-09, 1.227503e-07, -1.694195e-07, -5.592152e-08, 1.768714e-07, 
    -4.118328e-08, -2.495528e-08, -2.908837e-08, 6.527943e-09, 7.101589e-08, 
    -1.23822e-08, -4.065816e-08, -2.208708e-08, -4.992421e-08, -3.805053e-08, 
    4.383196e-09, -6.892492e-08, 5.254992e-08, 5.511106e-08, -7.921905e-09, 
    -1.819126e-08, -4.687836e-08, 1.817799e-08, -3.538349e-08, 1.38696e-07, 
    -6.697871e-08, 1.344434e-07, -1.078149e-09, -1.637488e-07, 4.315223e-08, 
    -3.619448e-09, 2.385377e-09, -9.091309e-08, 1.152728e-07, 2.758594e-08, 
    7.663061e-09, -3.414929e-08, -1.618758e-09, 5.9869e-08, -2.548119e-07, 
    -6.149987e-07, -1.765059e-08, 1.714704e-08, 3.94665e-08, -6.53253e-08, 
    1.250909e-07, -8.024621e-09, -6.533613e-08, 3.188212e-09, 3.982586e-08, 
    1.036585e-08, 5.419622e-08, -2.338766e-09, -4.306992e-08, -5.969014e-08, 
    -2.765637e-08, -9.894165e-09, -2.345473e-09, 3.900823e-09, 5.160359e-09, 
    6.199445e-09, 3.698844e-09, -1.450651e-09, -7.681678e-11, -3.00422e-08,
  1.988582e-08, 1.529431e-07, -6.214538e-08, -1.122288e-08, -8.990804e-08, 
    -9.612114e-08, -1.39126e-08, -2.862237e-09, 4.878001e-08, 7.980418e-09, 
    -1.218992e-07, -4.934697e-08, 2.490941e-08, 1.803522e-08, 3.417489e-08, 
    7.983005e-08, -3.892327e-08, 2.580072e-08, -1.946509e-08, -2.559449e-08, 
    1.915566e-09, -1.549267e-09, 3.885287e-08, -1.645009e-08, 8.562495e-09, 
    -9.498251e-09, 3.509268e-08, 9.750181e-09, -1.298317e-07, -5.401154e-08, 
    1.397183e-08, -1.068252e-07, -7.393277e-08, 2.383291e-08, -1.299856e-08, 
    -6.620161e-08, 2.017282e-08, 3.083755e-11, -1.827851e-08, -5.631679e-08, 
    1.09817e-07, 2.937992e-08, 1.723464e-09, 2.827329e-08, -3.268912e-08, 
    -1.178275e-07, -4.814922e-08, -4.229176e-08, -3.793249e-08, 4.251916e-09, 
    4.897146e-09, 6.653124e-09, 1.114183e-07, 2.871765e-08, -2.063226e-08, 
    -2.161187e-09, 9.188142e-08, -1.74615e-07, -6.462069e-08, 1.740439e-07, 
    -5.301894e-08, -2.441624e-08, 2.433296e-09, 4.306818e-08, 6.485674e-08, 
    -2.387054e-08, -7.915048e-09, -2.091764e-08, 8.504514e-09, -3.142981e-08, 
    1.126756e-08, -1.515758e-08, -1.52928e-07, -2.62213e-09, -9.285145e-09, 
    -3.358281e-08, -3.623195e-08, 1.488863e-08, -6.177972e-08, 1.879692e-07, 
    -5.167692e-08, 9.547476e-08, -2.174482e-08, 5.306475e-08, 2.004441e-08, 
    3.394365e-08, -1.609083e-07, -1.032731e-07, 1.185591e-07, 1.439554e-08, 
    1.226852e-09, -3.203044e-08, -7.642541e-09, 5.65975e-08, -2.78687e-07, 
    -6.195578e-07, -1.21585e-08, 2.74834e-08, 4.348811e-08, -4.459138e-08, 
    -1.368898e-08, -1.626545e-08, -8.716755e-08, -4.236966e-10, 7.105217e-08, 
    2.435064e-08, 6.508191e-08, 2.011234e-07, 1.252591e-07, -4.400277e-08, 
    -2.698965e-08, -8.99837e-09, 2.684885e-09, 3.417256e-09, 3.310276e-09, 
    4.712819e-09, 1.749981e-09, -9.180212e-10, -3.518892e-10, 1.393788e-07,
  -5.379616e-08, 2.477429e-08, -3.766809e-08, -1.715796e-08, 3.158789e-09, 
    -1.475382e-08, 2.149102e-08, 3.35516e-08, 3.358298e-08, 2.642435e-08, 
    -3.619448e-08, -3.743708e-09, 3.137893e-08, 2.251556e-08, 3.069647e-08, 
    6.842144e-08, -4.3556e-08, 4.34045e-09, 3.918717e-08, 4.726701e-08, 
    5.991637e-09, -2.226443e-09, 3.790967e-08, -2.09177e-08, 1.135106e-08, 
    -1.758781e-08, 1.260727e-07, 7.1268e-09, -1.317939e-07, -8.894392e-08, 
    4.281242e-08, -1.684004e-07, 1.199612e-08, 1.813498e-08, -2.963395e-08, 
    8.299708e-09, 2.913788e-08, 1.23174e-09, -1.157787e-09, -5.957331e-08, 
    1.207463e-07, 8.449751e-08, -2.098611e-08, 2.089771e-08, -8.212737e-10, 
    -9.388737e-08, -4.588338e-08, -4.574056e-08, -3.557636e-08, 5.199077e-09, 
    5.86104e-09, 2.018692e-08, 1.038842e-07, 2.560884e-08, -1.953525e-08, 
    -3.913271e-09, 6.99207e-08, -1.592749e-07, -6.950286e-08, 6.40963e-08, 
    -5.664299e-08, -2.677973e-08, 2.053821e-08, 7.754549e-08, 5.84017e-08, 
    7.284143e-09, 6.92728e-08, -2.845093e-08, 4.258482e-08, -4.01202e-08, 
    8.24366e-09, -1.719525e-08, -6.710366e-08, -2.977617e-08, -9.132584e-09, 
    -3.769105e-08, -3.755048e-09, 1.28839e-08, -8.159483e-08, -6.666187e-08, 
    -2.321156e-08, 7.455239e-08, -4.440972e-08, 5.919901e-09, 2.040576e-08, 
    2.992681e-08, -2.665058e-08, -9.824589e-09, 1.059832e-07, 2.14863e-08, 
    -1.069338e-09, -2.304687e-08, -5.968559e-09, 6.535535e-08, -2.018628e-07, 
    -5.331324e-07, -8.525285e-09, 4.430569e-08, 4.776075e-08, -4.193494e-08, 
    -1.705275e-07, -2.003028e-08, -5.479215e-08, -2.284757e-09, 1.621421e-07, 
    2.701927e-08, 8.55058e-08, 3.13534e-07, 2.232756e-07, 3.782498e-08, 
    -2.296474e-11, 3.911055e-09, 1.320927e-09, 2.813294e-09, 3.716877e-09, 
    5.81266e-09, 2.292026e-09, -1.96739e-09, -4.93678e-10, 1.224447e-07,
  -5.407963e-08, 3.835396e-09, -3.057238e-08, -1.710777e-08, 3.292456e-08, 
    6.926535e-08, 3.183294e-08, 3.700558e-08, 3.51651e-08, 4.497571e-08, 
    4.89041e-09, 3.347679e-09, 3.06805e-08, 2.579367e-08, 2.878704e-08, 
    5.241198e-08, -3.262518e-08, 1.288601e-08, 7.87411e-08, 7.579609e-08, 
    6.736343e-09, -2.595527e-09, 3.857525e-08, -2.354824e-08, 1.038535e-08, 
    -2.12172e-08, 1.146674e-07, -6.469776e-08, -3.467397e-08, -2.08791e-08, 
    1.597361e-07, 7.282608e-09, 1.695232e-07, -2.078167e-08, -3.722738e-08, 
    3.861879e-08, 3.479215e-08, 1.659274e-09, -3.704486e-10, -6.45917e-08, 
    1.373676e-07, 8.371416e-08, -3.273507e-08, 2.336386e-08, 1.246376e-07, 
    -9.571392e-08, -4.62876e-08, -3.801085e-08, -3.324141e-08, 5.666969e-09, 
    7.106152e-09, 2.699909e-08, 1.050767e-07, 2.337616e-08, -1.905e-08, 
    -2.414538e-09, 6.664146e-08, -1.452435e-07, -7.276213e-08, 9.311108e-08, 
    -6.051829e-08, -2.853352e-08, 3.002611e-08, 2.998198e-08, 4.8602e-08, 
    -2.134208e-07, 2.201642e-07, 8.99189e-09, 6.642387e-08, -1.157247e-08, 
    -7.662209e-09, -1.418977e-08, -1.310292e-08, -3.694112e-08, 
    -7.597713e-09, -6.964586e-08, 5.91298e-09, 1.398988e-08, -7.234913e-08, 
    -8.366061e-08, -1.506703e-08, 6.462911e-08, -5.363881e-08, 6.524999e-09, 
    2.040503e-08, 6.309205e-08, 6.112106e-08, -1.565496e-08, 9.438034e-08, 
    2.312999e-08, -2.921126e-09, -1.350323e-08, -6.188202e-09, 6.40253e-08, 
    -9.08629e-08, -4.454147e-07, -1.676232e-09, 1.19013e-07, 6.193983e-08, 
    9.188e-09, -8.695935e-08, -2.463751e-08, -3.512093e-08, -2.825132e-09, 
    -6.064681e-09, 1.922018e-08, 1.637854e-07, 1.715491e-07, 1.185833e-07, 
    9.297531e-08, 4.656482e-08, 1.284951e-08, 4.526441e-10, 2.697504e-09, 
    1.028371e-08, 2.887214e-09, 3.737256e-09, -1.189896e-09, 2.681659e-10, 
    1.23891e-07,
  -4.343644e-08, -3.894911e-09, -3.031266e-08, -1.838123e-08, 1.581475e-08, 
    2.980573e-08, 3.314472e-08, 2.30574e-08, 3.560672e-08, 4.521962e-08, 
    2.060835e-08, 2.421189e-08, 3.028993e-08, 2.59671e-08, 2.509978e-08, 
    3.745391e-08, -2.758386e-08, 2.966163e-08, 9.771287e-08, 2.652371e-08, 
    6.427058e-09, -7.904646e-10, 3.862749e-08, -2.526951e-08, 1.102785e-08, 
    -2.332115e-08, 1.33575e-07, 2.737102e-08, -5.704055e-08, 2.764386e-08, 
    1.125535e-07, 8.717325e-08, 2.239248e-07, -6.048026e-09, -4.393507e-08, 
    3.26371e-08, 3.995094e-08, 1.775703e-09, 1.148464e-09, -6.744163e-08, 
    1.430653e-07, 8.560494e-08, -3.730412e-08, 1.991341e-08, -4.51746e-08, 
    -1.001079e-07, -4.723313e-08, -4.188936e-08, -3.110197e-08, 6.042427e-09, 
    7.474426e-09, 2.981471e-08, 1.079817e-07, 2.361915e-08, -1.881117e-08, 
    2.986383e-09, 1.206712e-07, -1.433126e-07, -7.494467e-08, 8.00121e-08, 
    -6.325411e-08, -2.992351e-08, 3.520358e-08, 2.65532e-08, 3.590014e-08, 
    -7.955873e-08, 4.602839e-08, -3.799414e-09, 9.838539e-08, -2.965771e-08, 
    1.256683e-08, -1.037495e-08, -1.167621e-08, -3.829916e-08, -6.601191e-09, 
    -4.67378e-09, 6.48059e-09, 1.338634e-08, -7.416929e-08, -8.832978e-08, 
    -1.168303e-08, 5.873122e-08, -6.277799e-08, 4.758249e-09, 1.985177e-08, 
    7.038227e-08, 6.48771e-08, -1.619571e-08, 7.947095e-08, 2.253751e-08, 
    -4.62353e-09, -6.944015e-09, -5.918395e-09, 6.10618e-08, 2.61366e-10, 
    -3.745792e-07, -1.601152e-08, 4.012713e-08, 6.847654e-08, 1.315409e-08, 
    -1.536739e-08, -2.621714e-08, -3.549539e-08, -3.00718e-09, -4.766275e-08, 
    2.031493e-08, 5.395066e-07, 6.410187e-08, 1.065689e-08, 4.024605e-08, 
    5.276013e-08, 1.245883e-08, 2.011802e-09, 2.071374e-09, 2.250215e-08, 
    4.383458e-09, -3.030365e-09, -7.770815e-10, -2.568186e-10, 1.213741e-07,
  -2.98848e-08, -6.270909e-09, -2.859036e-08, -2.057021e-08, 1.218569e-08, 
    1.480959e-08, 2.933763e-08, 3.68255e-08, 3.547626e-08, 4.565828e-08, 
    2.637677e-08, 3.526731e-08, 2.68281e-08, 2.395478e-08, 2.151302e-08, 
    2.837365e-08, -2.051808e-08, 2.901783e-08, 1.054897e-07, 2.084772e-08, 
    5.523646e-09, -1.565638e-09, 3.806764e-08, -2.652968e-08, 1.323775e-08, 
    -2.463611e-08, 1.252834e-07, 9.369666e-08, -1.177963e-07, 1.843256e-08, 
    8.929993e-08, 6.076226e-08, 1.963525e-07, -1.869711e-08, -4.74185e-08, 
    2.994449e-08, 4.429527e-08, 1.635698e-09, 4.253576e-08, -7.115835e-08, 
    1.476642e-07, 8.748731e-08, -3.928517e-08, 6.2679e-09, 2.341295e-08, 
    -1.100847e-07, -4.903387e-08, -4.305508e-08, -2.79569e-08, 5.984546e-09, 
    7.702965e-09, 3.138786e-08, 1.089271e-07, 2.424991e-08, -1.876333e-08, 
    5.925074e-09, 1.764991e-07, -1.49501e-07, -7.639319e-08, 7.203823e-08, 
    -5.980695e-08, -3.022654e-08, 3.719839e-08, 2.770249e-08, 2.452049e-08, 
    -2.368682e-08, 1.174413e-08, 9.859662e-09, 9.383331e-08, -3.008239e-08, 
    1.139034e-08, -6.243852e-09, 1.910968e-08, -3.795088e-08, -6.644896e-09, 
    2.448417e-09, 9.45019e-09, 1.245121e-08, -7.47517e-08, -8.92e-08, 
    -3.198994e-08, 5.442724e-08, -6.925239e-08, 3.771049e-09, 1.899235e-08, 
    6.917099e-08, 7.366117e-08, -1.588995e-08, 6.727321e-08, 2.327494e-08, 
    -8.308859e-09, -4.556194e-09, -5.702589e-09, 5.845214e-08, 3.39233e-08, 
    -3.246278e-07, -2.378878e-08, -4.270504e-08, 7.154159e-08, 1.632503e-08, 
    -2.137125e-08, -2.655602e-08, -3.274081e-08, -3.523752e-09, 
    -5.888745e-08, 2.126586e-08, 2.114965e-07, 3.781571e-08, -2.048245e-08, 
    -1.675329e-08, 3.235306e-08, 1.498449e-09, 6.102084e-09, 1.076444e-09, 
    1.295444e-08, -5.535981e-10, -5.733227e-10, -1.289692e-09, -2.96339e-10, 
    1.189558e-07,
  -3.808918e-08, -2.207344e-09, -2.665183e-08, -2.409183e-08, 5.082484e-09, 
    1.614353e-10, 3.101013e-08, 3.228502e-08, 3.510763e-08, 4.549565e-08, 
    2.842648e-08, 3.984928e-08, 2.507318e-08, 2.211527e-08, 1.891431e-08, 
    2.997085e-08, -1.012577e-08, 2.964134e-08, 1.082634e-07, 1.360308e-08, 
    4.173899e-09, -3.901278e-09, 3.663263e-08, -2.753222e-08, 1.544686e-08, 
    -2.325964e-08, 1.366222e-07, 3.012337e-08, -1.258923e-07, -2.136676e-08, 
    9.271912e-08, 4.629464e-08, 1.971978e-07, -1.388366e-08, -4.934623e-08, 
    2.380034e-08, 4.667045e-08, 7.490542e-10, 7.620497e-08, -7.442088e-08, 
    1.449043e-07, 9.032829e-08, -4.000015e-08, 6.239048e-09, 3.364971e-08, 
    -1.179894e-07, -5.027925e-08, -4.110268e-08, -2.383395e-08, 8.815789e-09, 
    7.853117e-09, 3.217224e-08, 1.088451e-07, 2.470811e-08, -1.879322e-08, 
    -3.915488e-09, 1.604294e-07, -1.538918e-07, -7.796397e-08, 6.626169e-08, 
    -5.690572e-08, -3.015475e-08, 3.822402e-08, 2.950328e-08, 2.145066e-08, 
    1.438366e-09, 1.863054e-08, 1.167928e-08, 4.307753e-08, -2.872343e-08, 
    1.087983e-08, -8.426468e-09, 2.88062e-08, -3.701757e-08, -6.806403e-09, 
    7.525614e-09, 1.083424e-08, 1.171406e-08, -7.206283e-08, -8.857819e-08, 
    -3.049161e-08, 5.049719e-08, -7.390133e-08, 3.074547e-09, 1.703188e-08, 
    6.774758e-08, 7.958079e-08, -1.528497e-08, 5.627652e-08, 1.525098e-08, 
    -1.0863e-08, -2.592515e-09, -5.600555e-09, 5.613267e-08, 5.587663e-08, 
    -2.896331e-07, -3.177488e-08, -6.077357e-08, 7.439871e-08, 1.449416e-08, 
    -1.731451e-08, -2.704428e-08, -3.22656e-08, -6.33483e-09, -6.117602e-08, 
    2.193451e-08, -2.170132e-07, 2.444244e-08, -3.877904e-08, -2.994921e-08, 
    5.198899e-09, -1.463695e-08, 7.036078e-09, -4.42833e-09, 2.273737e-11, 
    2.53217e-09, 1.445841e-09, 1.065011e-09, -9.512178e-10, 1.167214e-07,
  -5.453012e-08, -1.94018e-09, -2.50551e-08, -2.744753e-08, 2.427441e-09, 
    -9.331984e-09, 3.279399e-08, 3.813261e-08, 3.317507e-08, 4.330082e-08, 
    2.88918e-08, 4.172591e-08, 2.547552e-08, 2.115269e-08, 1.959165e-08, 
    4.077819e-08, 1.56698e-09, 3.152667e-08, 1.086976e-07, 9.79162e-09, 
    2.157776e-09, -5.569063e-09, 3.417915e-08, -2.774402e-08, 1.653564e-08, 
    -2.209231e-08, 1.399324e-07, 2.906779e-08, -1.273238e-07, -2.31197e-08, 
    9.250596e-08, 4.359401e-08, 1.911542e-07, -1.431033e-08, -5.056211e-08, 
    1.641138e-08, 4.706372e-08, -1.060982e-09, 1.01048e-07, -7.24396e-08, 
    1.546511e-07, 9.330745e-08, -4.091419e-08, 9.558736e-10, 3.571688e-08, 
    -1.246686e-07, -5.160734e-08, -3.906055e-08, -2.045419e-08, 8.121951e-09, 
    7.275958e-09, 3.219952e-08, 1.09583e-07, 3.47404e-08, -1.888684e-08, 
    -3.650939e-09, 1.208576e-07, -1.579524e-07, -7.97132e-08, 6.768811e-08, 
    -5.528591e-08, -2.911338e-08, 3.885043e-08, 3.502851e-08, 1.502012e-08, 
    4.26644e-09, 3.375612e-08, 2.097761e-08, 2.9999e-08, -2.700654e-08, 
    1.067133e-08, 1.130252e-08, 3.593152e-08, -3.563957e-08, -7.133245e-09, 
    1.162834e-08, 1.111724e-08, 1.147814e-08, -5.608149e-08, -8.745496e-08, 
    -2.898469e-08, 4.682949e-08, -7.710867e-08, 2.50111e-09, 1.635715e-08, 
    6.64096e-08, 8.258269e-08, -1.417618e-08, 4.744059e-08, -2.353488e-09, 
    -1.060926e-08, -2.38772e-09, -5.679738e-09, 5.231011e-08, 7.438246e-08, 
    -2.615254e-07, -3.312116e-08, -7.321273e-08, 7.390747e-08, 1.450469e-08, 
    -1.431135e-08, -2.717844e-08, -3.699021e-08, -5.800153e-09, 
    -6.179323e-08, 2.292779e-08, -2.173624e-07, 1.84657e-08, -4.934031e-08, 
    -3.574735e-08, -2.582738e-09, -2.267564e-08, 3.491436e-09, -1.177057e-08, 
    -5.38796e-09, -1.004753e-09, 3.469438e-10, -6.805596e-09, -1.366011e-09, 
    1.143922e-07,
  -6.622031e-08, -1.373564e-09, -2.288061e-08, -3.219418e-08, -3.293508e-10, 
    -1.413798e-08, 3.292996e-08, 4.208539e-08, 3.130151e-08, 4.145943e-08, 
    2.734828e-08, 4.205015e-08, 2.537399e-08, 1.905232e-08, 1.959802e-08, 
    -3.849351e-09, 1.340156e-08, 3.189984e-08, 1.069976e-07, 6.647269e-09, 
    -1.336389e-09, -7.879862e-09, 3.018783e-08, -2.726995e-08, 1.712806e-08, 
    -2.067804e-08, 1.384237e-07, 2.739353e-08, -1.273214e-07, -2.455999e-08, 
    9.319933e-08, 4.39702e-08, 1.892729e-07, -1.967476e-08, -5.105755e-08, 
    1.023079e-08, 4.666635e-08, -4.36728e-10, 2.449094e-07, -6.66819e-08, 
    1.524494e-07, 9.47465e-08, -4.206623e-08, -1.527848e-09, 3.460673e-08, 
    -1.327163e-07, -5.310659e-08, -3.557122e-08, -1.865819e-08, 7.474249e-09, 
    5.558505e-09, 3.129389e-08, 1.112168e-07, 2.396009e-08, -1.903599e-08, 
    -1.427338e-10, 7.930055e-08, -1.563169e-07, -8.159599e-08, 6.805126e-08, 
    -5.273e-08, -2.739478e-08, 3.823061e-08, 3.916069e-08, 2.358433e-09, 
    5.312586e-09, 4.341882e-08, 1.894102e-08, 1.640615e-08, -2.487275e-08, 
    1.011745e-08, 6.973175e-08, 4.153435e-08, -3.338107e-08, -7.622113e-09, 
    9.159635e-09, 1.097742e-08, 1.075131e-08, -5.558234e-08, -8.439372e-08, 
    -2.910713e-08, 4.318255e-08, -7.385751e-08, 1.750891e-09, 1.668343e-08, 
    6.511084e-08, 8.673157e-08, -1.226226e-08, 4.025256e-08, -3.379404e-08, 
    -1.111687e-08, -2.941897e-09, -5.768641e-09, 4.852049e-08, 8.850861e-08, 
    -2.275972e-07, -3.462824e-08, -7.666927e-08, 7.39002e-08, 1.397746e-08, 
    -1.10914e-08, -2.775695e-08, -3.575204e-08, -5.488772e-09, -6.093626e-08, 
    2.438753e-08, -2.125362e-07, 1.636295e-08, -5.519212e-08, -3.776961e-08, 
    -6.225264e-09, -2.450668e-08, -3.228251e-09, -1.773765e-08, 
    -7.117364e-09, 9.766268e-10, -8.437311e-09, 3.628351e-10, -3.315414e-09, 
    1.111728e-07,
  -7.321199e-08, -1.155911e-09, -2.120686e-08, -3.966323e-08, -6.149492e-09, 
    -1.861002e-08, 3.039742e-08, 4.113559e-08, 2.901794e-08, 3.844167e-08, 
    2.4332e-08, 4.034706e-08, 2.192752e-08, 1.432437e-08, 1.745963e-08, 
    -3.969166e-08, -1.609284e-08, 2.991459e-08, 1.016135e-07, 5.800587e-09, 
    -6.942116e-09, -1.307529e-08, 2.152848e-08, -2.745531e-08, 1.736504e-08, 
    -1.817938e-08, 1.490624e-07, 2.451208e-08, -1.213543e-07, -2.760629e-08, 
    9.694446e-08, 4.169175e-08, 1.871588e-07, -3.234226e-08, -5.022815e-08, 
    3.313573e-09, 4.601605e-08, -9.309247e-10, 4.067393e-07, -5.444375e-08, 
    1.752122e-07, 9.289312e-08, -4.166066e-08, -2.745608e-09, 2.940175e-08, 
    -1.351452e-07, -5.441876e-08, -3.135915e-08, -1.843517e-08, 4.423157e-09, 
    1.39292e-09, 2.815733e-08, 1.143436e-07, 2.551884e-08, -1.930296e-08, 
    2.996842e-09, 5.006706e-08, -1.593534e-07, -8.283388e-08, 6.424264e-08, 
    -4.747261e-08, -2.439646e-08, 3.450879e-08, 3.904698e-08, -5.305045e-08, 
    4.328342e-09, 3.76229e-08, 1.869063e-08, 1.71313e-08, -2.650444e-08, 
    8.654581e-09, 1.035081e-07, 3.448901e-08, -2.885207e-08, -8.416318e-09, 
    -1.985194e-08, 1.061153e-08, 9.919859e-09, -4.837685e-08, -7.675629e-08, 
    -2.888947e-08, 3.875831e-08, -7.586669e-08, 3.688569e-10, 1.356904e-08, 
    6.269153e-08, 7.438308e-08, -7.967344e-09, 3.538439e-08, -1.041691e-07, 
    -1.383245e-08, -2.981404e-09, -6.044161e-09, 4.276279e-08, 9.943284e-08, 
    -1.786602e-07, -3.457311e-08, -7.89077e-08, 7.216346e-08, 1.382738e-08, 
    -6.01284e-09, -2.902758e-08, -3.153046e-08, -5.071897e-09, -5.696319e-08, 
    2.743701e-08, -2.011238e-07, 1.797008e-08, -5.767714e-08, -3.697295e-08, 
    -7.534879e-09, -2.530436e-08, -4.487163e-09, -2.196629e-08, 
    -8.362065e-09, 5.20447e-10, -8.769774e-09, 3.251728e-10, -8.654979e-09, 
    1.046181e-07,
  -3.813435e-13, 1.318128e-14, 3.127335e-13, 3.832741e-13, 2.816013e-13, 
    2.580164e-13, 4.995097e-13, 4.208786e-13, 2.066691e-14, -4.199629e-13, 
    -3.466237e-13, 6.421277e-13, 1.926948e-14, -9.412352e-15, -5.944987e-14, 
    1.927168e-13, -4.131467e-13, -4.59323e-13, -1.740986e-14, -2.790713e-14, 
    -1.330227e-12, -1.898941e-12, -2.1436e-13, 4.434029e-13, -6.268589e-13, 
    -1.670106e-14, 7.661897e-14, 2.881742e-15, -5.193835e-14, -7.639518e-14, 
    8.663629e-14, 7.927895e-14, -1.805262e-14, -6.097799e-14, 3.055864e-14, 
    -1.169428e-13, 2.502757e-13, -3.972646e-12, -4.748487e-13, -1.352254e-13, 
    1.031201e-13, -4.832435e-13, 1.439434e-13, 4.706655e-14, 1.726154e-13, 
    4.128777e-14, 4.333976e-13, 3.493857e-13, 1.742305e-12, 1.009577e-12, 
    -2.099032e-12, -1.488581e-13, -4.794843e-13, -2.573653e-13, 
    -1.219653e-13, -1.568955e-12, -3.674547e-13, 5.365039e-13, 2.318162e-13, 
    1.817704e-13, 1.041513e-12, 2.176464e-14, 5.708961e-13, -2.922166e-12, 
    -2.136336e-12, 2.054921e-13, -4.362359e-14, -5.479449e-15, 1.708511e-13, 
    1.149659e-13, -2.60706e-14, 1.163244e-13, 1.323816e-13, -3.526638e-14, 
    5.399249e-13, 2.16398e-14, 3.777345e-14, -1.688334e-12, -1.4525e-12, 
    -5.535135e-13, -6.676394e-14, -1.658024e-12, 1.653889e-12, -4.652386e-13, 
    3.675449e-13, 4.735891e-14, 1.223629e-13, -1.575043e-13, -5.29361e-13, 
    -3.371995e-13, 6.853029e-13, 1.810989e-12, 1.142479e-12, -1.247465e-14, 
    1.00034e-13, 4.300427e-13, 3.905135e-13, 5.720969e-13, 2.468971e-13, 
    2.152628e-13, -1.563694e-12, 1.757091e-13, -1.848668e-12, 5.417673e-13, 
    -1.284739e-13, 2.013838e-13, -5.695553e-14, -2.398165e-13, -2.747589e-13, 
    -6.311224e-14, -7.193561e-14, -7.223389e-14, 5.539523e-14, -4.567752e-14, 
    6.953307e-13, -1.663511e-12, 1.963763e-12, -2.899043e-13, 3.725126e-13, 
    -1.68591e-12,
  1.180844e-13, 2.71404e-14, -7.871146e-14, -1.553856e-13, -9.028058e-14, 
    -1.404769e-14, 6.624071e-14, 2.135499e-13, 1.105138e-13, 1.368168e-13, 
    1.797349e-13, -1.634236e-13, 1.556771e-13, -1.243214e-13, -1.271279e-13, 
    6.769806e-14, -1.230505e-13, -5.018838e-14, -1.432143e-13, -2.000631e-13, 
    -3.498106e-13, -1.185e-12, -6.783114e-13, 3.000819e-13, -3.373725e-14, 
    -2.914413e-13, -8.688574e-13, -1.466172e-13, -6.777158e-14, 
    -1.610734e-13, 5.466476e-14, 2.326024e-13, -2.89216e-14, 2.103259e-15, 
    4.781908e-14, -1.058701e-13, -1.572336e-13, 4.741472e-14, 1.857014e-13, 
    3.56455e-13, -8.174148e-13, 2.538752e-13, -1.644945e-13, 3.131364e-14, 
    -1.20756e-12, -2.372742e-12, -9.429873e-13, -2.224939e-14, -5.378726e-13, 
    2.46765e-13, 8.128986e-14, 5.773336e-14, -2.721772e-13, -2.478028e-12, 
    2.986279e-14, -1.383619e-12, -1.222883e-13, -1.215675e-12, -3.874949e-13, 
    -2.590228e-12, 3.884475e-13, -1.332706e-13, -4.002764e-14, -3.818942e-14, 
    -8.100739e-14, 4.440943e-13, 2.580031e-14, 1.452109e-14, -1.360599e-13, 
    1.696889e-13, -2.019766e-13, 1.664162e-13, 1.252547e-13, -9.905533e-14, 
    1.541778e-12, -3.684091e-13, -1.293724e-13, 5.433777e-13, 1.638725e-12, 
    -1.017054e-12, -3.212898e-13, 6.663214e-13, -1.68685e-12, 3.344571e-14, 
    -6.49555e-13, -9.82294e-13, -7.353201e-13, 4.743879e-13, 3.880301e-14, 
    -3.564699e-13, 1.335362e-13, 4.129636e-13, 5.62945e-13, -9.743735e-13, 
    1.10656e-13, 9.251665e-13, -9.50969e-14, -1.803256e-13, 4.092433e-13, 
    -5.187524e-13, 2.926553e-13, -4.754449e-13, -3.607491e-13, -2.504309e-12, 
    2.446708e-13, 7.104718e-13, 2.456569e-13, 1.135833e-12, 4.018665e-13, 
    -1.569803e-15, -1.30413e-13, -1.579914e-13, -1.16528e-13, -5.134971e-14, 
    -1.505162e-13, -6.303351e-13, -5.49028e-13, 5.352965e-12, -2.161446e-13, 
    -5.590455e-15,
  5.479645e-14, -9.153095e-14, -1.820349e-13, -1.638689e-13, 2.997602e-15, 
    1.780451e-13, 3.49748e-13, 3.261488e-13, 2.269643e-13, 4.361095e-14, 
    -5.647566e-14, -5.07927e-14, 1.415534e-15, 2.102485e-14, 7.920054e-14, 
    -4.696868e-14, -1.787417e-13, -2.173019e-13, -3.448561e-13, -2.06779e-14, 
    8.011716e-13, 5.775311e-13, 4.129752e-13, 3.180095e-14, 3.750264e-13, 
    9.810833e-13, 3.642781e-13, 1.63744e-13, 1.142003e-13, 1.68969e-13, 
    3.394507e-14, -5.134781e-15, -9.554857e-15, -1.022793e-14, 3.180789e-14, 
    1.793496e-13, -2.728571e-12, 3.787014e-13, -1.487976e-13, 6.75477e-13, 
    2.079836e-13, -1.440084e-12, -2.513042e-13, 9.516975e-14, -1.500328e-13, 
    5.578871e-13, -5.414211e-13, 1.038912e-12, -3.065534e-13, -6.984387e-14, 
    3.685238e-13, -3.796546e-13, 1.974385e-12, -2.242066e-11, 5.594483e-14, 
    -1.2336e-12, -2.41758e-13, -1.162271e-12, 7.612299e-13, -4.751781e-13, 
    1.236039e-12, -8.901352e-13, 1.229711e-13, -1.822445e-13, -1.746214e-13, 
    -1.70565e-13, 3.700651e-13, 4.760081e-14, -5.515727e-14, 5.12923e-14, 
    -8.596526e-13, 8.434919e-14, 1.025915e-12, 1.136868e-13, -5.598848e-13, 
    4.874781e-13, -1.527077e-13, 8.787415e-13, -4.3988e-12, -9.780926e-13, 
    1.074339e-12, 5.294883e-13, 1.018949e-12, 5.156292e-13, -1.738193e-13, 
    6.774928e-13, 2.918568e-13, 2.735798e-13, -3.626008e-13, 9.243648e-13, 
    -1.552994e-13, -2.162645e-13, 4.304005e-13, -1.173489e-12, -2.730455e-14, 
    -4.134068e-13, -5.216689e-13, -1.644518e-13, 6.06272e-13, 1.578471e-12, 
    -7.753867e-13, 2.46195e-13, 5.159796e-13, 2.501341e-13, -2.043851e-13, 
    -4.567804e-13, -4.319461e-13, -7.160592e-13, -1.141275e-12, 
    -1.997152e-12, -1.450014e-12, -4.513473e-13, -3.66214e-13, -1.306108e-13, 
    -6.983789e-13, -9.376646e-13, -7.623841e-12, 1.62623e-11, -1.06513e-12, 
    3.15685e-13,
  8.061607e-14, 1.180028e-13, 8.174017e-14, 1.261213e-13, 2.69243e-13, 
    3.870931e-13, 4.189843e-13, 2.391698e-13, -1.181832e-13, -4.392736e-13, 
    -2.115391e-13, -4.894279e-13, -4.230366e-13, -8.444911e-13, 
    -8.778672e-13, -3.324896e-13, -5.239975e-14, -6.503825e-14, -3.41371e-13, 
    -3.347045e-13, -1.146583e-13, -2.867151e-14, 1.427192e-13, -3.307771e-13, 
    -1.327216e-12, -1.703762e-12, -6.419865e-14, 1.791761e-13, 3.552436e-13, 
    4.566347e-13, -1.055822e-13, -1.539463e-13, -1.107323e-12, -2.32897e-13, 
    -1.273287e-13, -9.010848e-14, -2.039914e-12, 1.111937e-12, 1.857403e-13, 
    1.712991e-13, 4.672374e-14, 1.515857e-12, -4.307145e-13, -1.392656e-13, 
    2.140094e-13, -2.88658e-14, -1.299599e-12, 4.354607e-13, 8.54411e-13, 
    1.123421e-12, -4.128798e-13, 4.182765e-13, 2.013417e-13, 2.755923e-12, 
    2.477782e-13, 6.108725e-13, -1.912748e-12, -6.082399e-13, 1.87797e-13, 
    1.096817e-12, 3.448908e-13, 3.100298e-14, -8.331391e-13, -1.394357e-13, 
    -2.020328e-13, 2.903511e-13, -2.424588e-13, -3.711892e-13, -4.957146e-14, 
    -2.440131e-13, -1.236788e-13, 3.27488e-13, -2.134959e-13, 3.622658e-13, 
    -9.889714e-13, 6.203787e-13, 2.095176e-12, 2.234945e-12, -2.368588e-11, 
    3.513856e-14, 1.189278e-12, -4.826799e-14, -1.677686e-13, -2.299591e-12, 
    -4.25715e-13, -4.722195e-13, -4.899275e-13, -9.826862e-14, -1.977815e-13, 
    -3.184883e-13, -1.508932e-13, -1.759381e-12, 7.428537e-13, -3.776188e-13, 
    -2.164519e-13, -4.477546e-12, -1.085451e-12, 1.122019e-13, -7.638418e-12, 
    -2.803796e-12, 4.223427e-13, -1.857924e-12, 5.991024e-13, 2.507794e-13, 
    -4.364703e-13, -1.822847e-13, -3.113482e-13, -4.527073e-13, 
    -2.619294e-13, -6.785544e-13, -6.208367e-13, -4.909823e-13, 
    -1.805361e-13, 8.962275e-14, -8.965051e-15, 5.373701e-13, 4.314065e-12, 
    1.338377e-12, -6.563847e-14, -9.964529e-13,
  8.365114e-13, 5.114381e-13, 4.141826e-13, 4.037187e-13, 3.986672e-13, 
    4.26173e-13, 7.654571e-13, 9.218321e-13, 6.959572e-13, -9.505868e-13, 
    -6.071671e-13, -7.017303e-13, -8.314183e-14, -2.865763e-14, 7.687601e-13, 
    -2.278122e-13, -4.327871e-13, -6.264433e-13, -2.865173e-13, 
    -4.187345e-13, -1.505879e-13, -7.533557e-13, -1.14149e-12, -1.004571e-12, 
    -1.785086e-12, -1.467701e-12, 1.119868e-12, 4.283379e-13, 8.507084e-15, 
    8.13058e-13, 8.086448e-13, 6.022544e-13, 1.188077e-13, -7.345374e-13, 
    -8.923556e-13, -4.97255e-13, -9.871632e-13, 1.573977e-12, 6.674244e-13, 
    -2.338518e-13, -3.215123e-13, 2.272488e-13, -4.103315e-13, -2.40051e-13, 
    5.099671e-13, 5.079964e-13, 2.299549e-14, -1.721394e-12, 1.246545e-12, 
    1.641288e-11, 9.721043e-14, 1.518161e-12, -2.575801e-13, -1.458492e-12, 
    1.90252e-13, 1.716405e-13, 2.950126e-12, -1.682549e-12, -1.01158e-13, 
    2.217879e-13, -1.6806e-14, -4.703044e-13, -2.117057e-13, -4.588025e-13, 
    -6.497608e-13, 1.918882e-13, -1.506156e-13, 1.146999e-13, 4.331396e-13, 
    -1.360315e-12, 4.407447e-13, -3.993056e-13, -4.869022e-13, -2.175898e-13, 
    -2.087663e-13, 5.551809e-13, 2.406686e-13, -5.700232e-13, -7.078481e-12, 
    3.149564e-13, 1.08788e-13, 5.723644e-13, -3.765321e-13, -1.787001e-12, 
    -9.563322e-13, -1.271899e-13, 1.06512e-13, 1.195294e-13, -5.001065e-13, 
    1.050729e-12, -2.968598e-13, 2.032055e-12, 4.935705e-13, 1.601372e-12, 
    -4.300588e-13, 1.235709e-11, -3.430173e-13, -2.808725e-13, -2.65489e-12, 
    -1.433437e-13, 3.067976e-12, 6.431487e-13, 1.594117e-12, 1.486415e-13, 
    -3.307493e-13, -4.162642e-13, -2.451234e-13, 1.696282e-13, -5.237616e-13, 
    -5.183215e-13, -1.819517e-13, 2.840922e-13, -8.59729e-14, 1.752348e-13, 
    7.495393e-14, 2.002537e-12, 9.71628e-12, -1.295723e-11, -1.244014e-12, 
    -6.259299e-13,
  8.576473e-14, 1.647571e-13, 1.511846e-13, 1.656175e-13, 5.009604e-13, 
    4.97935e-13, 6.305789e-13, -1.326717e-14, -8.049117e-16, -1.135203e-14, 
    -1.224021e-14, -7.155387e-14, -1.553119e-12, -3.022027e-12, 
    -7.422118e-13, -5.489525e-13, -2.242267e-12, -3.302636e-13, 
    -8.213048e-13, -1.396716e-12, -2.016248e-12, -8.577306e-13, 
    -1.647543e-12, -1.717571e-12, -2.19863e-12, -2.231881e-12, -1.905115e-12, 
    -5.269118e-13, -6.016854e-13, -1.980777e-12, -3.4375e-12, -2.761569e-12, 
    -1.998041e-12, 1.131484e-12, -1.938893e-12, 4.71817e-13, -6.06043e-13, 
    1.776357e-13, 1.398132e-12, 2.606498e-13, 1.489037e-12, -2.201656e-12, 
    -1.027123e-12, -8.73402e-13, 8.442691e-12, 8.753276e-13, -4.116707e-13, 
    2.18936e-13, -6.765366e-13, 8.365558e-12, -2.529921e-13, -2.074979e-12, 
    3.107514e-13, 9.139856e-13, 3.128234e-13, -2.591954e-13, -8.679168e-14, 
    1.005807e-13, 3.895023e-13, -4.060398e-13, -2.041228e-12, -2.681466e-12, 
    5.575262e-13, -2.559975e-12, -1.920097e-12, -4.949652e-13, 7.418788e-13, 
    3.519074e-12, 7.634088e-12, 1.532829e-12, 1.65043e-12, -6.414036e-13, 
    -1.051104e-13, -2.439715e-13, -5.750231e-12, -6.017409e-14, 
    -5.589487e-13, -3.522183e-14, -1.942777e-12, 2.276374e-12, 1.474071e-12, 
    5.374125e-13, 1.720013e-13, -1.347616e-12, 1.652567e-13, -3.260142e-12, 
    -8.200385e-13, -1.704192e-14, 6.386805e-13, -1.684305e-12, -2.840506e-13, 
    -3.13638e-14, -5.04527e-14, 2.692888e-12, 4.118372e-13, -1.762784e-13, 
    -2.107536e-13, -1.545153e-13, 1.278391e-11, 6.631529e-13, 1.419698e-12, 
    -1.365895e-12, 1.43041e-12, -1.200449e-12, -2.380318e-13, -4.313216e-13, 
    -1.331213e-12, -1.43302e-13, -4.401479e-13, -3.283485e-13, 1.887379e-14, 
    1.651179e-13, 5.966061e-13, 2.122191e-12, -7.053247e-13, 2.47101e-12, 
    2.739468e-12, -2.033405e-12, -1.611732e-13, -3.535228e-13,
  -1.133316e-12, -9.611756e-13, 7.577272e-14, -1.823541e-13, 5.532796e-13, 
    4.847234e-13, -1.59317e-14, 1.001199e-12, 7.382983e-14, -6.126211e-12, 
    -7.933487e-12, -1.032019e-11, -5.546286e-12, -9.830303e-12, 
    -4.764522e-12, -1.944506e-12, -5.845269e-13, -1.015965e-12, 
    -1.475001e-12, -2.484901e-12, -2.149725e-12, -1.216194e-12, 9.220402e-14, 
    1.259326e-12, 4.662937e-14, -2.01561e-13, -5.67818e-12, -4.970468e-12, 
    7.301382e-13, -9.699908e-12, -1.497191e-12, 2.614131e-12, -3.436307e-12, 
    3.372302e-12, 1.384781e-12, 4.764189e-12, -1.105804e-12, -1.956768e-15, 
    -5.967449e-14, -1.509826e-12, 2.908118e-13, 1.072031e-12, -1.618247e-12, 
    -6.167072e-13, 4.164835e-12, 6.288359e-12, 2.997325e-13, 1.821265e-12, 
    1.24708e-12, -6.380854e-12, 2.942702e-12, -1.881773e-12, 2.558143e-12, 
    8.923762e-12, -1.030898e-13, 2.770006e-13, -3.586187e-12, -2.025491e-13, 
    1.628841e-12, -1.197951e-12, 2.394474e-12, -5.346334e-12, -5.234702e-13, 
    -2.118528e-12, -3.105516e-13, 1.516537e-11, 1.448519e-11, -8.627543e-13, 
    -2.776945e-12, 1.43352e-12, 1.720513e-12, -2.820577e-12, -2.159661e-12, 
    -4.95437e-13, -4.379769e-12, -4.924949e-13, -4.938758e-13, -7.619738e-13, 
    -9.399321e-12, -4.528988e-12, 4.738404e-12, 4.373034e-12, 1.012301e-12, 
    -2.771672e-13, 3.651801e-12, -1.021283e-11, 4.48086e-12, -6.583623e-13, 
    -8.077514e-13, -4.352907e-13, -4.993284e-12, -2.388045e-12, 
    -8.856804e-14, 8.774592e-13, 2.21595e-12, 5.970335e-13, 1.512612e-12, 
    -2.053357e-13, 1.835199e-11, 3.126677e-12, 1.614819e-13, 4.954023e-13, 
    3.875372e-14, -6.385014e-12, -1.382228e-13, 7.972512e-13, 2.396972e-13, 
    1.69631e-12, 2.059464e-13, -7.101542e-13, 3.587131e-13, 3.169742e-12, 
    1.316613e-12, 2.534084e-13, 3.204048e-12, 1.064099e-12, 1.100071e-12, 
    8.528612e-13, -6.791408e-13, -3.654077e-12,
  -2.063127e-12, 3.842981e-12, 8.861467e-12, 1.080275e-11, 1.171108e-11, 
    9.27225e-12, 1.116052e-11, 4.922174e-13, -1.671052e-12, 6.94883e-12, 
    -1.261286e-11, -2.44752e-11, -1.017003e-11, -1.528766e-11, -1.278327e-11, 
    2.097528e-12, 3.025413e-13, -7.948642e-12, 1.508321e-12, -7.502887e-13, 
    -6.508682e-13, -3.594347e-13, 2.445266e-13, -2.743361e-13, 1.697087e-12, 
    1.43166e-11, 1.668526e-11, -1.442735e-13, 1.866174e-12, 2.736311e-12, 
    3.223977e-12, -1.077455e-11, -4.367673e-12, -4.220346e-12, 6.892431e-12, 
    1.034856e-11, -5.467143e-12, -4.705403e-13, -2.118716e-11, 5.374923e-13, 
    4.890843e-12, -2.342626e-12, -8.5848e-13, -1.623338e-12, 1.745382e-12, 
    6.721568e-12, 1.545986e-12, -4.236889e-13, 3.682144e-12, -1.083391e-11, 
    3.885503e-13, -4.491074e-12, -8.384071e-13, 7.690504e-12, -4.261161e-13, 
    4.645728e-13, 7.735979e-12, 6.948498e-13, 2.136935e-12, 1.188218e-11, 
    -2.270073e-11, 9.037215e-13, -6.458722e-13, 5.866974e-13, -3.824286e-12, 
    4.854611e-11, 1.339956e-11, 8.50664e-12, 8.174295e-12, 1.650524e-11, 
    -3.816114e-12, 1.342332e-11, 1.699252e-12, -5.879186e-13, -4.578948e-13, 
    -1.603717e-13, -4.415357e-13, 8.373857e-14, -1.554484e-11, -1.383904e-11, 
    1.003517e-11, -2.649866e-11, 2.912892e-12, 1.442674e-11, 1.382783e-13, 
    -7.904621e-12, 7.493672e-12, 2.085609e-12, -1.092659e-13, 8.965884e-13, 
    -1.723732e-12, -8.676804e-12, 1.916939e-13, 5.14766e-13, 4.843514e-12, 
    -1.374434e-12, 3.637668e-12, -3.301803e-13, 1.606548e-12, -2.880807e-13, 
    7.668255e-12, 1.65e-12, -5.753523e-13, -4.057586e-11, -5.305201e-13, 
    1.492306e-12, 2.986111e-12, 1.632749e-12, 4.456435e-13, 1.203593e-12, 
    6.143752e-12, 2.156719e-12, -4.652945e-12, -7.95175e-12, -3.256839e-12, 
    -1.304062e-12, 9.510726e-13, -2.862807e-12, -2.596881e-14, 2.04875e-12,
  2.340572e-12, 9.099221e-12, 1.905159e-11, 1.973871e-11, 1.422301e-11, 
    5.515755e-12, 1.07237e-11, 3.770467e-11, 2.619144e-11, 4.199141e-12, 
    4.989065e-12, -1.912082e-12, -1.00786e-12, 3.221978e-12, -8.690881e-12, 
    2.058204e-12, -3.489747e-12, -1.564554e-12, 7.349538e-13, -1.248557e-12, 
    -2.528644e-12, 1.059153e-13, 3.695932e-12, -7.310874e-12, 5.155321e-13, 
    9.530432e-12, 3.324452e-12, 4.385159e-12, -2.732981e-12, 9.614531e-12, 
    8.245071e-13, -7.929213e-12, 2.306766e-12, -4.209022e-12, -5.331124e-12, 
    1.66589e-12, -9.485967e-13, -8.201426e-13, 1.883171e-11, 1.95538e-12, 
    -1.575906e-12, -6.687095e-12, 2.582795e-13, 5.064677e-12, 7.425505e-12, 
    2.725542e-12, 2.146894e-13, -7.11764e-13, -7.230882e-14, -6.428854e-12, 
    -4.857503e-13, 1.731948e-12, 1.599054e-13, 3.065326e-14, -1.341141e-12, 
    1.490474e-13, 5.976053e-12, 1.522132e-12, -1.601635e-12, 1.448766e-11, 
    -5.058892e-11, 2.914224e-12, 7.049361e-13, -4.681e-12, -8.301981e-12, 
    9.470646e-12, -4.28213e-13, 7.336964e-12, -2.645123e-11, 2.344791e-13, 
    2.702283e-13, 7.756684e-12, 5.508649e-12, -5.906109e-12, 3.78007e-12, 
    2.274292e-13, -3.036668e-13, 1.703471e-12, -1.194979e-11, 1.263378e-12, 
    5.203782e-12, 1.286833e-11, 1.270956e-12, -2.909339e-11, -9.836076e-12, 
    -3.095968e-12, 1.004025e-11, 7.255863e-13, 6.906229e-13, -7.671641e-14, 
    -8.881562e-12, -1.274678e-11, 1.456474e-13, 1.670758e-12, -2.338019e-12, 
    3.653078e-12, -1.981304e-12, -1.381023e-11, -4.60848e-12, -1.601175e-12, 
    2.545131e-12, -2.054308e-12, 7.515343e-13, -4.600983e-11, 2.239653e-12, 
    6.052381e-13, 6.519008e-12, 3.285316e-12, 1.574019e-12, 1.197653e-12, 
    -2.167988e-12, -1.455197e-11, 7.840228e-12, 1.694805e-11, -1.727468e-11, 
    -8.483492e-13, 1.422334e-13, -1.644429e-12, 4.918808e-13, 7.812362e-12,
  -1.580458e-12, 6.918799e-12, 9.857726e-12, 6.573686e-12, 7.47935e-12, 
    3.589995e-11, 2.119638e-11, -2.354084e-11, 3.383005e-11, -8.005985e-12, 
    -5.356826e-14, 8.78736e-12, -4.347606e-11, -3.984174e-11, -3.476219e-12, 
    -3.480438e-13, -6.911721e-12, -4.598127e-12, 7.937748e-13, 3.385625e-12, 
    -1.932843e-12, 7.082002e-12, 1.746203e-11, 1.26682e-12, 8.27044e-12, 
    -9.876933e-12, -3.889666e-12, -2.895623e-11, -5.317691e-12, 1.147077e-11, 
    1.120931e-11, 2.644224e-11, 7.485401e-12, 2.21399e-11, -3.560957e-11, 
    3.52437e-11, 3.334338e-12, -7.404077e-13, 1.56089e-11, 8.10274e-13, 
    5.909162e-12, 6.453893e-12, 7.936485e-12, 7.342215e-12, 7.424339e-12, 
    -2.142347e-11, -4.645728e-13, -1.064884e-12, -9.304113e-12, 3.997924e-12, 
    6.49758e-14, 6.392831e-12, 2.882217e-12, -2.997824e-13, -2.555338e-12, 
    5.295209e-13, 5.846101e-12, 3.061496e-13, -2.227196e-12, 4.244674e-12, 
    -4.123968e-11, 3.335388e-12, -2.717937e-12, -6.3484e-12, -4.777678e-12, 
    -2.320366e-14, 2.234407e-11, -2.624534e-11, -3.069134e-11, 1.040217e-10, 
    -1.37611e-11, -9.333118e-11, 1.21308e-11, 3.438527e-12, -4.064138e-13, 
    8.826273e-15, -4.139467e-13, 1.245865e-12, -7.189901e-13, -5.540013e-12, 
    5.906109e-13, 4.080048e-11, -2.662037e-13, -2.374712e-11, 1.047273e-12, 
    -3.625322e-12, -1.313727e-12, 8.102186e-12, 5.366029e-13, -3.188477e-12, 
    -1.061945e-11, -4.797595e-12, -1.469797e-13, 4.609041e-12, -1.18423e-11, 
    -4.936163e-13, -2.837286e-12, 4.086342e-12, -1.917982e-11, -2.993317e-12, 
    -2.159373e-11, -6.995297e-12, -4.174612e-13, -2.678378e-11, 
    -9.812096e-12, 1.088629e-12, 8.255063e-13, -2.909728e-12, 1.593892e-12, 
    -3.960887e-12, -8.724299e-12, -1.377065e-11, 3.879508e-11, 1.664247e-11, 
    -1.398776e-11, -6.680434e-13, -3.166911e-14, -2.552389e-12, 4.274327e-12, 
    1.093736e-12,
  1.995848e-12, 5.737633e-12, 1.307732e-12, 7.946677e-11, 2.6534e-11, 
    4.302303e-11, -4.619638e-13, -2.351674e-11, 2.504996e-12, 2.056222e-11, 
    -1.51168e-12, -1.149603e-11, -1.019296e-11, -4.473777e-11, -1.765543e-11, 
    -1.643041e-12, -6.23871e-12, -2.974065e-12, 6.398312e-12, 3.383849e-12, 
    7.377432e-13, -1.053091e-11, 5.81768e-12, -1.43574e-11, -4.349743e-12, 
    6.23831e-11, -8.614254e-11, 1.385458e-11, -9.596768e-13, -2.691103e-11, 
    1.893186e-11, 2.578382e-11, 8.306689e-12, 2.295253e-11, 3.383183e-12, 
    3.392187e-11, -2.759681e-13, -5.469097e-13, -1.629041e-11, -3.83249e-13, 
    1.552505e-11, 1.675649e-11, 2.27468e-12, 1.98337e-12, 9.218182e-13, 
    -2.534961e-11, -6.403766e-13, -2.43508e-12, -4.997158e-12, 1.52877e-12, 
    4.415052e-12, -2.992473e-11, 3.648359e-12, -7.800427e-14, -2.452621e-13, 
    5.164758e-13, -4.520828e-13, -2.612799e-13, -3.834377e-13, -8.339732e-12, 
    -1.751943e-11, -3.874678e-12, 2.595812e-12, -4.844835e-12, -4.64595e-12, 
    2.56728e-12, 2.798406e-11, -6.858025e-11, -9.901413e-11, -2.658185e-11, 
    -2.67959e-11, 8.189116e-11, 1.426814e-11, 1.510514e-11, -3.431355e-12, 
    -5.462297e-13, -3.784334e-13, -4.696529e-11, 2.495296e-12, 1.245781e-12, 
    -2.582656e-12, 1.311328e-11, -9.851564e-13, -4.513723e-12, -4.830469e-12, 
    -1.496069e-10, 2.191247e-11, 1.445521e-11, -1.190693e-12, -5.842105e-12, 
    -2.597877e-11, -9.072432e-12, 1.292577e-13, -2.534282e-11, -3.024359e-12, 
    2.412737e-13, -6.042433e-12, -6.023015e-11, -1.928524e-11, -3.446865e-12, 
    -1.67335e-11, -8.874387e-12, -1.584149e-12, -6.197487e-12, -1.335587e-11, 
    -3.849365e-12, -4.735656e-12, -1.624623e-11, -1.81688e-12, -8.280265e-12, 
    -1.712019e-11, -6.981526e-12, 2.595968e-11, 1.896416e-11, 2.855494e-13, 
    -1.451728e-13, -2.071954e-14, -2.291264e-12, 9.131557e-12, -2.195355e-12,
  -9.679813e-12, 6.18553e-11, 6.099965e-11, 4.504142e-11, 5.712431e-12, 
    -1.699418e-11, -2.030687e-11, -4.187417e-11, -1.359313e-10, -4.4169e-11, 
    -5.194456e-11, 5.017831e-11, -1.384348e-11, 8.31446e-13, -9.524048e-12, 
    -1.74728e-12, -4.468448e-12, -2.852107e-12, -5.277723e-14, 9.528822e-12, 
    7.775558e-12, -1.605127e-11, 2.134681e-11, 1.188716e-12, 1.370905e-10, 
    1.532374e-11, -8.828727e-11, -3.040213e-11, -5.414003e-12, -4.755785e-11, 
    -3.240874e-11, 2.595701e-11, 9.178081e-11, -6.139755e-12, -2.939338e-11, 
    5.648604e-11, -1.815481e-12, -3.590461e-13, 2.099532e-11, -4.118705e-13, 
    1.158087e-11, 5.542566e-12, 8.540196e-12, 3.792505e-13, 4.663647e-11, 
    8.630319e-12, -1.497358e-12, -4.047485e-12, 9.098389e-12, 5.18266e-14, 
    1.31589e-11, -5.325029e-11, 2.97381e-12, 4.231726e-13, 1.538769e-13, 
    5.92304e-14, 7.330359e-12, -5.880186e-13, -2.579981e-12, 8.729087e-12, 
    -3.214318e-12, -3.758771e-12, -3.477441e-12, -3.571188e-12, 
    -2.546563e-12, -5.578205e-12, 7.375345e-11, -1.506505e-10, -5.310863e-12, 
    -4.239631e-11, -2.017275e-13, 7.805145e-11, -3.368406e-11, 1.027789e-11, 
    -5.277245e-12, -7.293055e-13, -2.373796e-13, -3.020098e-11, 5.664191e-13, 
    4.287681e-12, -6.339873e-12, -8.964051e-13, 1.527445e-12, -4.13517e-11, 
    -1.780531e-11, -8.601431e-11, 4.322731e-11, 2.437128e-11, -4.16155e-12, 
    -5.114797e-13, -2.308376e-11, -2.16207e-12, 1.489198e-12, -4.3565e-11, 
    1.590872e-11, 2.265599e-12, -7.778823e-12, 1.963962e-11, -2.763267e-11, 
    -3.8195e-12, 1.673084e-11, 3.181365e-12, -2.201274e-12, 8.168952e-13, 
    1.497757e-11, -3.369971e-12, -3.736711e-11, -3.80691e-11, -1.52649e-11, 
    -2.087885e-11, -2.393441e-11, -3.483658e-12, 1.467926e-11, 3.706846e-11, 
    1.599998e-11, 4.583001e-14, 1.133676e-13, -7.413757e-13, 5.072484e-12, 
    -3.326395e-11,
  8.772316e-12, 7.373213e-11, 2.17022e-11, -2.172618e-11, -4.191647e-11, 
    -3.31537e-11, -3.020895e-11, -1.76545e-10, -2.922835e-10, -3.04037e-10, 
    7.247314e-12, 1.47486e-10, -8.194734e-11, -1.015898e-11, -1.813816e-11, 
    -1.235212e-12, -6.628898e-12, -7.86593e-12, 1.185996e-13, 2.468914e-11, 
    5.448975e-12, -1.150813e-11, 5.829714e-11, -1.399769e-12, 2.484124e-10, 
    -1.382983e-11, -1.229434e-10, -4.483125e-11, -4.765766e-11, 
    -7.156542e-11, -3.448775e-11, 5.013256e-11, 1.325311e-10, -3.991607e-11, 
    -1.707043e-10, -1.482126e-11, 3.37308e-13, -1.98952e-13, 4.459477e-11, 
    1.40199e-13, 2.672173e-12, 1.170553e-11, 1.695871e-11, -2.696142e-13, 
    1.091824e-10, 4.747891e-11, -2.417733e-12, -2.604306e-12, 4.170575e-12, 
    2.064043e-13, 2.969369e-11, -4.56053e-11, 1.69198e-12, 1.060707e-12, 
    1.495915e-13, -4.971579e-13, 7.677192e-11, -4.920508e-13, -6.814061e-12, 
    1.843437e-11, -6.189937e-12, 1.550493e-11, -5.098366e-12, -5.043788e-12, 
    -7.323031e-12, -1.177529e-10, 1.231009e-10, -4.127365e-11, -2.61251e-11, 
    -7.300827e-13, -5.268008e-12, 8.512013e-11, 4.827916e-12, 3.061063e-11, 
    -6.065148e-12, -2.406964e-13, -1.701417e-13, -1.471745e-11, 
    -1.249889e-13, -2.301492e-12, -9.747092e-12, -1.708145e-12, 2.553957e-12, 
    -1.177074e-10, -7.282064e-11, -5.977041e-11, 1.023384e-10, 3.04663e-11, 
    -2.184621e-12, 3.489764e-12, -3.188916e-11, 2.336797e-13, 1.973643e-12, 
    -1.664196e-11, 2.007772e-11, -2.717382e-13, -6.358913e-12, 5.130318e-11, 
    -4.28293e-11, -3.085798e-12, 4.589107e-11, 2.273778e-11, -2.219433e-12, 
    5.155598e-13, 1.557643e-11, 2.279998e-11, -5.483658e-11, -5.651724e-11, 
    -2.071188e-11, -1.818234e-11, -2.775469e-11, -6.424639e-12, 2.379008e-11, 
    5.137046e-11, 1.897105e-11, -1.240119e-13, 3.41116e-13, 3.866699e-13, 
    1.719236e-12, -4.232859e-11,
  5.742606e-11, -1.899236e-11, -3.282175e-11, -2.30207e-11, 5.325518e-12, 
    -3.79563e-11, -8.759082e-11, -2.562013e-10, -7.271339e-11, -2.942402e-11, 
    1.365263e-11, 8.515988e-11, -1.250844e-10, -2.791722e-11, -2.986056e-12, 
    -8.951062e-13, -9.503909e-12, -7.621459e-12, 2.495576e-11, 2.631806e-11, 
    5.025758e-12, 1.289102e-11, 3.827871e-11, -1.236744e-11, 1.682672e-10, 
    2.584435e-10, -1.714899e-10, -3.785727e-11, -9.951373e-11, -3.996359e-11, 
    -1.024199e-10, 9.483614e-11, 1.052993e-10, 1.66529e-11, -1.096794e-10, 
    -2.862417e-10, 2.921219e-13, -1.948997e-13, -2.223328e-10, 2.513634e-12, 
    -5.656009e-12, 2.994405e-11, 1.237643e-11, -1.729172e-13, 1.359286e-10, 
    -3.117062e-11, -2.056133e-13, -6.883383e-13, 1.268319e-12, -9.367507e-14, 
    4.969625e-11, -5.385381e-11, -3.925749e-13, 4.469225e-12, 3.78364e-13, 
    -1.361133e-13, -7.633494e-11, -4.805934e-13, -2.21374e-12, 9.755474e-12, 
    -1.64242e-11, 7.951462e-11, -2.696066e-11, -8.422241e-12, -7.927436e-12, 
    -7.712995e-10, 8.552448e-11, -2.0556e-11, 2.074252e-11, 5.5973e-12, 
    -5.632694e-11, 8.624346e-11, 1.908083e-10, 7.544587e-11, -3.97824e-12, 
    2.522427e-13, -1.34337e-14, -2.148925e-11, -1.057732e-12, 5.374901e-11, 
    -1.078115e-11, 1.86704e-12, 4.094503e-13, -1.147589e-10, -1.744067e-10, 
    -2.621396e-10, 1.033782e-10, 3.485656e-11, -3.842343e-13, -2.879919e-13, 
    -1.333555e-11, 7.249579e-12, 1.31839e-12, -1.376321e-12, 1.003375e-11, 
    -8.101297e-12, -4.527934e-13, 6.534417e-11, -2.673506e-11, -2.655032e-12, 
    9.116796e-11, 6.489415e-11, -1.863815e-12, 7.68996e-13, -3.685496e-11, 
    5.012346e-11, 6.219913e-12, -7.984591e-11, -2.283462e-11, -4.591882e-12, 
    -2.931078e-11, -9.73488e-12, 4.271694e-11, 4.56053e-11, 1.263967e-11, 
    -7.953638e-14, 8.789636e-13, 1.958989e-13, 5.539735e-13, -8.721912e-12,
  5.670442e-11, -5.697842e-11, 1.582379e-11, 9.030554e-11, -2.036593e-12, 
    -9.680479e-11, -1.201808e-10, -2.709064e-10, -1.364868e-10, 
    -5.560885e-11, -2.222844e-11, 2.40945e-11, 1.378848e-10, -4.802958e-11, 
    4.323697e-11, -3.213429e-13, -9.815171e-12, 9.894308e-13, 3.362038e-11, 
    2.675371e-11, -7.647216e-13, 5.66005e-11, -5.780665e-11, -1.086158e-10, 
    1.48666e-10, 1.828564e-10, -1.924731e-10, -4.299849e-11, -6.959278e-11, 
    -6.33662e-11, -1.108624e-10, 8.413847e-11, 6.483702e-11, 2.419647e-10, 
    1.409819e-10, -2.461906e-10, 5.328627e-13, -2.326472e-13, -4.647487e-10, 
    8.428947e-12, -2.398863e-11, 4.530287e-11, 1.505185e-11, -3.700582e-13, 
    2.561e-10, -5.1398e-11, 3.830936e-12, 3.410827e-12, 4.736655e-13, 
    -8.296697e-13, 5.780032e-11, -5.073675e-11, -1.175371e-12, 4.49667e-12, 
    4.691026e-13, 4.154455e-13, 4.230336e-10, -9.80993e-14, -1.67546e-12, 
    -1.90446e-11, -2.411671e-11, 1.590315e-10, -7.223866e-11, -7.528467e-12, 
    1.495959e-12, 5.226766e-10, 3.58483e-10, -6.238698e-11, 6.395373e-11, 
    2.759615e-11, -1.5608e-10, 3.387246e-11, 3.997473e-10, 1.351763e-10, 
    -9.488499e-12, 1.193268e-12, 1.140754e-13, -1.435496e-11, -3.863132e-13, 
    1.205325e-10, -1.009792e-11, 7.211531e-12, -2.006395e-12, -1.436042e-10, 
    -2.334177e-11, -6.841954e-10, -1.514158e-10, 4.35616e-11, -1.79351e-12, 
    -4.657386e-12, -1.446265e-11, 1.225384e-11, 5.759837e-13, -1.059286e-11, 
    -2.030953e-11, -2.136331e-11, 7.452705e-12, 7.611511e-11, -3.901324e-12, 
    4.072298e-13, 1.409814e-10, 7.945386e-11, -1.114248e-12, 6.576684e-13, 
    -4.795142e-11, -3.748557e-11, 5.988854e-11, 5.996981e-12, -1.982947e-11, 
    7.568612e-12, -2.544498e-11, -4.584333e-12, 5.833245e-11, 2.267342e-11, 
    3.579359e-12, -1.005418e-13, 1.634082e-12, -7.979728e-14, 2.249589e-13, 
    1.642726e-10,
  4.271294e-11, -2.233458e-11, 1.306799e-10, 8.681011e-11, -2.982281e-11, 
    -2.718137e-11, -7.688739e-11, -2.954628e-10, -3.211773e-10, 
    -3.380767e-10, -2.545764e-10, 2.215388e-10, 9.647763e-10, -5.645218e-11, 
    8.928724e-11, 8.593126e-13, -6.84226e-12, 1.072564e-11, 2.502165e-11, 
    4.332668e-11, -5.858869e-12, 6.191447e-11, -2.157647e-10, -2.930087e-10, 
    6.869594e-10, 1.154333e-09, -9.956036e-12, -7.5564e-11, -3.247047e-11, 
    -1.024749e-10, -1.385527e-10, -2.847034e-10, 1.439697e-10, -7.165712e-10, 
    2.623364e-10, -7.190715e-10, 1.937117e-12, -2.484679e-13, -6.848935e-10, 
    2.154286e-11, -8.724212e-11, 4.479217e-11, 3.94853e-11, -6.197584e-12, 
    3.845728e-10, -4.052625e-11, 1.045342e-11, 3.64142e-11, -5.775025e-12, 
    -2.495004e-12, 4.170597e-11, -6.182566e-11, 2.438938e-12, -1.077867e-11, 
    1.464606e-13, -7.371881e-14, 9.274701e-10, -1.23368e-13, -3.284599e-11, 
    -6.430712e-11, -2.886624e-11, 1.878768e-10, -6.232659e-11, 6.816769e-13, 
    1.520446e-11, -9.445555e-11, 2.262204e-10, -1.632072e-11, 2.867706e-11, 
    2.972067e-11, -1.917857e-10, -6.145795e-11, 2.632157e-10, 1.143836e-10, 
    -2.344533e-11, 1.981082e-12, 7.605028e-14, -5.700551e-12, 4.180034e-12, 
    1.918674e-10, -1.457412e-11, 9.750844e-12, -4.823697e-12, -1.454405e-10, 
    6.339951e-11, -7.611729e-10, -6.230083e-11, 5.772316e-11, -4.318837e-12, 
    -3.610445e-13, 6.184786e-11, -6.146292e-11, 3.723688e-13, -2.149099e-11, 
    -5.452838e-11, -4.568097e-11, 1.801661e-11, 1.360911e-11, -1.380673e-12, 
    4.14202e-12, 1.371965e-10, 1.392122e-10, -3.724243e-13, 4.652945e-13, 
    2.087619e-11, 6.541878e-12, 3.945155e-11, 1.67296e-10, -7.092549e-12, 
    7.295942e-12, -1.399725e-11, 7.079226e-12, 6.903944e-11, 1.973222e-11, 
    -7.256862e-12, -1.230127e-13, 2.44349e-12, 2.908229e-13, -1.472378e-12, 
    3.136793e-10,
  3.180811e-11, 1.484746e-11, 1.045393e-10, 1.104332e-10, 1.837435e-10, 
    1.869871e-10, -3.641643e-11, -3.733842e-10, -1.634846e-10, -4.195553e-10, 
    -2.387186e-10, 8.890655e-10, 8.846583e-10, -7.555845e-11, -4.877454e-11, 
    4.218981e-12, -5.49294e-13, 1.7782e-11, 1.792677e-11, 6.18694e-11, 
    -1.20306e-11, 4.491763e-11, -2.729117e-10, -3.352565e-10, 1.420054e-09, 
    2.094176e-09, 1.140232e-10, -1.159848e-10, 4.119662e-10, -1.869502e-10, 
    -2.646516e-10, -3.414364e-10, 4.031508e-11, -4.938738e-11, 3.561282e-10, 
    -1.277745e-09, 3.878986e-12, 4.152234e-14, -1.157852e-09, 5.753438e-11, 
    -3.100763e-10, 2.949352e-11, 7.78797e-11, -1.748718e-11, -3.565082e-11, 
    -2.622642e-10, 1.865419e-11, 1.493021e-10, -2.647416e-11, -4.091838e-12, 
    3.763612e-11, -1.038913e-10, 1.651563e-11, -3.568563e-11, 3.648015e-12, 
    -3.936851e-13, 9.482786e-10, -2.338441e-12, -1.212703e-10, -1.169671e-10, 
    -3.706835e-11, 1.751956e-10, 1.169087e-11, 7.521761e-12, 2.00195e-11, 
    -1.087159e-10, 3.566096e-10, 1.529354e-11, 2.137934e-11, -1.374656e-11, 
    -1.066838e-10, -3.756573e-11, 1.873637e-10, -5.623702e-11, -5.252834e-11, 
    1.489253e-12, 6.972201e-14, 6.623591e-13, 1.058487e-11, 2.767642e-10, 
    -3.459122e-11, 1.709646e-11, -5.420775e-12, -3.45451e-10, 9.307288e-11, 
    6.690892e-11, -5.948242e-11, 7.231971e-11, 8.429368e-13, 3.252576e-11, 
    2.725347e-10, -9.972898e-11, -1.088019e-14, -2.475091e-11, 4.498335e-11, 
    -7.775794e-11, 1.111888e-11, 5.357736e-11, 6.383782e-13, 5.446621e-12, 
    1.157356e-10, 2.640959e-10, 3.459455e-13, 2.565836e-12, 1.81799e-11, 
    1.029778e-10, -1.968232e-10, -1.939988e-10, -1.202356e-10, 9.587664e-12, 
    5.164535e-12, 1.562372e-11, 6.850054e-11, 3.976441e-11, -2.295164e-11, 
    8.204548e-13, 3.47633e-12, 1.379064e-12, -4.647283e-12, 3.292182e-10,
  6.932765e-11, 9.046097e-11, 1.524345e-10, 3.551115e-11, 1.636931e-10, 
    4.845173e-10, 2.583871e-10, -5.66196e-10, 3.12177e-11, 9.77245e-11, 
    1.049898e-09, 1.133794e-09, -1.761327e-09, -1.500613e-10, -1.069882e-10, 
    9.85576e-12, 1.094911e-11, 2.055156e-11, 1.682809e-11, 7.49143e-11, 
    -1.851497e-11, 3.722533e-11, -2.532214e-10, -2.329159e-10, 1.807416e-09, 
    2.451317e-09, 1.054747e-10, 1.92788e-11, 1.364922e-09, -2.661711e-10, 
    -7.332552e-10, -6.279119e-10, -2.768026e-10, -7.602843e-10, 2.940919e-10, 
    -1.818096e-09, -2.934897e-12, 2.427392e-12, -1.717881e-09, 1.455623e-10, 
    -5.99665e-10, -1.889688e-11, 1.064908e-10, -2.575759e-11, 4.745324e-10, 
    -6.090684e-10, 2.437428e-11, 3.482188e-10, -5.960282e-11, -7.050915e-12, 
    1.716556e-10, 1.516831e-11, 4.557528e-11, -3.963905e-11, 2.409397e-11, 
    -1.154632e-12, 7.969518e-10, -2.202149e-12, -2.630633e-10, -1.990528e-10, 
    -5.422329e-11, 1.373799e-10, 3.201528e-11, 8.911982e-12, 2.167617e-11, 
    2.771898e-10, 2.502157e-09, 5.934755e-10, 9.299761e-11, -9.928591e-11, 
    -4.728129e-11, -2.825473e-11, 6.614478e-10, -3.65814e-10, -1.009402e-10, 
    -1.096012e-12, 5.386802e-13, 4.009237e-12, 1.419447e-11, 3.807372e-10, 
    -7.607603e-11, 5.645373e-11, -2.16005e-12, -5.868923e-10, -2.004938e-10, 
    1.494213e-09, -2.160174e-10, 8.778578e-11, 3.923489e-11, 7.366374e-11, 
    2.042366e-10, -7.210801e-11, -2.317702e-12, -6.215917e-11, 1.72065e-10, 
    -9.683898e-11, -2.055849e-11, 2.542695e-10, -4.447998e-12, 5.892886e-12, 
    -3.049472e-11, 3.943057e-10, 1.093126e-12, 1.25755e-11, -1.988294e-10, 
    1.732676e-10, -3.031655e-10, -1.001419e-09, -4.869989e-10, 3.003287e-11, 
    2.664535e-11, 1.42375e-11, 7.467449e-11, 1.220766e-10, -9.867662e-12, 
    3.525891e-12, 3.799183e-12, 3.221201e-12, -6.038947e-12, 2.664375e-10,
  2.475247e-10, 2.841105e-10, 3.588454e-10, 7.641177e-11, -1.514131e-10, 
    1.559393e-10, 8.179732e-10, -6.045155e-10, 2.374634e-11, 2.066507e-10, 
    1.724427e-09, -1.309321e-09, -2.079808e-09, -2.946337e-10, -1.427622e-10, 
    7.198153e-12, 2.754632e-11, 1.846523e-11, 9.506618e-12, 6.982859e-11, 
    -2.728129e-11, 4.957101e-11, -2.464908e-10, -6.158736e-10, 1.892616e-09, 
    3.573184e-09, -8.576251e-11, -3.444853e-10, 4.22844e-10, -5.017888e-10, 
    -1.669648e-09, -3.701928e-12, -8.983498e-10, -9.875905e-10, 1.355076e-10, 
    -2.75989e-09, -2.551879e-11, 7.583267e-12, 4.229506e-10, 3.246921e-10, 
    -7.638611e-10, -7.581846e-11, 1.197513e-10, -2.907297e-11, 6.417054e-10, 
    -1.288651e-09, 2.702016e-11, 5.213163e-10, -8.890808e-11, -1.461964e-11, 
    3.03447e-10, 4.426539e-10, 8.824124e-11, -5.732232e-11, 5.592114e-11, 
    -3.039347e-12, -6.776695e-10, 8.430234e-12, -3.177164e-10, 1.749547e-10, 
    -9.050538e-11, 9.15783e-11, 1.750884e-10, 9.474377e-12, 2.479297e-11, 
    1.700521e-09, -2.318949e-09, 1.078558e-09, 3.046097e-11, -2.094964e-10, 
    -2.694165e-10, 8.021708e-10, 9.522445e-10, -7.393801e-10, -7.602417e-11, 
    -4.455103e-12, 2.18936e-12, 1.348788e-11, 1.77188e-11, 5.7614e-10, 
    -1.063754e-10, 1.010474e-10, 3.751666e-12, -5.301324e-10, -4.877556e-10, 
    1.596383e-09, -2.372502e-10, 1.04432e-10, 1.075359e-10, 1.232436e-11, 
    2.804512e-11, -6.398295e-11, -7.156942e-12, -1.322313e-10, 7.550724e-10, 
    -8.614016e-11, -7.663346e-11, 5.511929e-10, -2.08118e-11, 6.974688e-12, 
    -2.32852e-10, 4.245466e-10, -1.462608e-12, 3.365819e-11, -6.45219e-10, 
    1.034337e-10, 4.495355e-10, -8.607977e-10, -4.105516e-10, 2.004157e-10, 
    4.688516e-11, 1.216804e-11, 1.094129e-10, 2.258318e-10, 3.143441e-11, 
    6.580692e-12, 4.678924e-12, 4.792056e-12, -5.735856e-12, 1.820801e-10,
  3.160636e-10, 4.11724e-10, 5.214176e-10, 2.582681e-10, 2.472333e-10, 
    -3.453096e-10, 9.145111e-10, -5.328147e-10, -8.684964e-11, -7.459917e-10, 
    5.788863e-10, -1.430465e-10, -4.321876e-10, -4.051799e-10, -2.379963e-10, 
    -3.002754e-11, 3.242633e-11, 1.05409e-11, -9.461765e-12, 6.61089e-11, 
    -4.467182e-11, 2.985701e-11, -2.068532e-10, -2.131415e-09, 1.955364e-09, 
    5.648182e-09, 1.604832e-10, -1.613991e-09, -5.857075e-10, -7.170726e-10, 
    -2.740975e-09, 5.559357e-10, -1.520014e-09, -1.547271e-09, 2.823626e-10, 
    -2.595172e-09, -8.019185e-12, 1.437339e-11, 4.795417e-09, 6.547424e-10, 
    -3.432732e-10, -6.438938e-11, 1.423555e-10, -3.375911e-11, -2.618634e-10, 
    -1.766182e-09, 5.771739e-11, 5.249117e-10, -8.497949e-11, -2.874989e-11, 
    2.008385e-10, 1.565468e-10, 6.787744e-11, -5.683915e-11, 6.240289e-11, 
    -5.968559e-12, -1.689301e-09, 2.815099e-11, 5.236699e-12, 3.786464e-10, 
    -1.518714e-10, 4.445155e-11, 1.97744e-10, 6.264145e-12, 2.740847e-11, 
    3.28712e-09, -2.51012e-09, 1.535383e-09, -1.20837e-09, -4.019967e-10, 
    -7.666969e-10, 1.264652e-09, 1.367873e-09, -9.04457e-10, 8.19604e-11, 
    -6.65068e-12, 5.946355e-12, 3.05036e-11, 3.584368e-11, 7.522587e-10, 
    -8.639134e-11, 1.582132e-10, 8.586909e-12, -4.470522e-10, -2.2753e-10, 
    6.772964e-10, 2.332001e-10, 1.184546e-10, 8.634593e-11, -2.183391e-10, 
    1.035119e-10, -5.583303e-11, -1.39444e-11, -5.902479e-11, 2.125468e-09, 
    -6.757191e-11, -1.546056e-10, 6.603997e-10, -2.615508e-11, 9.126211e-12, 
    -2.776233e-10, 3.023621e-10, -1.051115e-11, 6.060841e-11, -1.113982e-09, 
    -4.319318e-10, 7.079919e-10, -1.140769e-09, -2.144688e-09, 9.06283e-10, 
    9.289636e-11, 1.363532e-11, 5.953638e-11, 2.561649e-10, 7.572964e-11, 
    1.041869e-11, 1.06759e-11, 4.776401e-12, -2.743583e-12, 1.121592e-10,
  -6.068035e-12, 1.143661e-09, 1.07211e-09, -7.135412e-10, 3.34353e-10, 
    5.745591e-10, -3.040412e-10, 3.042402e-10, -2.045795e-10, -1.251408e-09, 
    4.284431e-10, -5.798313e-10, 2.15195e-10, -3.936265e-10, -4.181118e-10, 
    -2.887987e-10, -5.967706e-11, 5.044853e-12, 1.494804e-11, 7.075585e-11, 
    -6.711787e-11, -3.791456e-11, -1.439844e-10, -2.279208e-09, 2.748308e-09, 
    3.778894e-09, 4.46434e-10, -3.62121e-09, 5.613288e-11, -7.251799e-11, 
    -4.634316e-09, 1.720011e-09, -2.028912e-09, -4.775544e-09, 4.833538e-10, 
    -1.901967e-09, 9.247287e-11, 1.723244e-11, 8.553315e-09, 1.155395e-09, 
    -1.240665e-10, 7.118217e-11, 1.996305e-10, -6.709544e-11, -9.591474e-10, 
    -1.722427e-09, 1.49619e-10, 3.537721e-10, -7.346444e-11, -6.596945e-11, 
    2.834373e-10, -2.534364e-10, -1.656929e-10, 2.707736e-11, 5.36911e-11, 
    -8.412826e-12, 5.559656e-09, 4.420144e-11, 8.485515e-10, 2.160476e-10, 
    -2.240341e-10, -6.197354e-11, 3.518608e-11, 2.751221e-12, 1.983551e-11, 
    3.044789e-09, -9.364953e-12, 3.24674e-09, -3.059995e-09, -7.800907e-10, 
    -1.745477e-09, 6.170751e-09, -2.221725e-10, -1.148919e-09, 7.85505e-11, 
    -8.000711e-12, 1.261036e-11, 1.250875e-10, 5.843184e-11, 1.946034e-10, 
    -2.196998e-11, 3.149989e-10, 1.315925e-11, -5.677663e-10, 2.155218e-10, 
    -1.031992e-09, 5.641994e-10, 1.137153e-10, -1.802973e-10, -4.770655e-10, 
    2.65743e-10, -3.113882e-11, -1.569944e-11, 3.821157e-11, 1.558135e-09, 
    -7.80787e-11, -2.148852e-10, 4.149854e-10, 2.359002e-12, 1.24885e-11, 
    -3.073382e-10, 1.434319e-10, -2.433609e-11, 8.94298e-11, -1.151108e-09, 
    -1.387548e-09, -1.012353e-09, 2.826965e-10, 2.143992e-10, 1.538012e-09, 
    1.153495e-10, -7.099743e-11, 9.507062e-12, 3.278444e-11, 7.212009e-11, 
    1.703313e-11, 2.251355e-11, 3.229417e-12, 4.973799e-13, 2.576428e-11,
  -4.690648e-10, 3.142794e-09, 1.053095e-10, -3.836355e-09, -4.586902e-09, 
    6.850698e-10, -1.11104e-09, 1.234106e-09, 3.776535e-11, -1.80286e-10, 
    1.382567e-09, -6.622756e-10, 4.750902e-10, -3.234888e-10, -7.048229e-10, 
    -7.604655e-10, -1.019984e-10, 6.536993e-12, 9.134382e-11, 1.320544e-10, 
    -9.890044e-11, -1.16934e-10, -3.274891e-11, -3.814691e-10, 4.367472e-09, 
    -1.620442e-09, 4.309875e-09, -6.309584e-09, -9.40048e-12, 2.116352e-10, 
    -6.290826e-09, 1.571387e-09, -1.115133e-09, -9.729249e-10, 3.47093e-10, 
    -4.750227e-09, 2.816705e-10, 1.948308e-11, 6.779821e-09, 1.470566e-09, 
    -3.956686e-10, 1.564828e-10, 2.341345e-10, -3.12431e-10, -7.639969e-10, 
    -1.028546e-09, 2.146834e-10, 2.698712e-10, -2.194966e-10, -8.178169e-11, 
    4.276117e-10, -5.092957e-10, -5.15719e-10, 2.969998e-10, 1.256073e-10, 
    -6.210144e-12, 1.011956e-08, 4.39087e-11, 1.715674e-09, -3.064944e-10, 
    -1.777849e-10, -1.878604e-10, 3.969802e-11, 3.602451e-12, -5.765344e-12, 
    3.319094e-09, 1.29738e-10, 3.028156e-09, -2.850335e-09, -1.376399e-09, 
    -9.42471e-10, 1.173793e-08, 5.457679e-11, -1.166704e-09, 8.149357e-11, 
    2.110312e-12, 2.234657e-11, 3.973817e-10, 4.522711e-11, -3.037073e-10, 
    5.068301e-11, 3.573884e-10, 2.529532e-11, 4.026006e-10, -7.556409e-10, 
    -1.563784e-09, 2.580762e-10, 9.232082e-11, -6.265033e-10, 7.045742e-11, 
    7.055689e-12, -2.250815e-10, -2.181366e-11, 7.284911e-11, 2.424805e-09, 
    -1.503878e-10, -2.530001e-10, 3.388649e-10, 5.095302e-11, 6.352252e-13, 
    -9.266685e-10, 2.24273e-10, -3.482548e-11, 1.269571e-10, -1.006008e-09, 
    -2.336101e-09, -2.337522e-09, -1.798313e-10, -2.599521e-10, 2.57473e-09, 
    2.939444e-10, -2.538982e-10, 6.222223e-11, 1.590905e-11, -5.591971e-12, 
    2.470841e-11, 5.540812e-11, 1.052936e-12, -5.214496e-12, -6.333067e-11,
  -1.008814e-09, 3.338783e-09, 2.596579e-09, 1.543029e-09, -9.149446e-09, 
    -6.889081e-09, 1.642249e-09, 1.142851e-09, 1.597826e-09, 2.127706e-09, 
    2.380546e-09, 2.367614e-09, 1.018392e-09, -3.000764e-10, -9.118253e-10, 
    -1.443823e-10, -4.324278e-10, 2.927436e-11, 1.331628e-10, 3.105356e-10, 
    -1.471108e-10, -1.896154e-10, 1.197691e-10, 5.254321e-10, 1.234241e-09, 
    -6.617483e-09, 8.365561e-09, -1.05391e-08, 1.489099e-09, 7.575565e-09, 
    -6.459061e-09, -1.243919e-09, 1.379689e-09, 8.005117e-10, 3.443432e-10, 
    -2.605745e-09, 3.955762e-10, 2.197709e-11, 2.86478e-09, 1.113018e-09, 
    -1.222037e-09, -9.210055e-11, 7.026983e-10, -5.349623e-10, 1.052925e-09, 
    -5.730527e-10, 1.856719e-10, 7.678551e-10, -6.4434e-10, -7.900525e-11, 
    4.23837e-10, -7.665335e-10, -7.56431e-10, 4.720107e-10, 4.442839e-10, 
    2.273737e-12, 3.721098e-09, 2.905267e-11, 2.456183e-09, -9.939303e-10, 
    -1.666223e-10, -2.420819e-10, 4.845901e-12, 8.599841e-11, -2.871729e-11, 
    5.653945e-09, -1.505214e-10, 2.712738e-09, -2.9587e-09, -1.79692e-09, 
    2.236931e-10, 1.389016e-08, 3.449259e-10, -9.495267e-10, 9.330535e-10, 
    2.292211e-11, 3.117506e-11, 8.335768e-10, 2.340279e-11, -8.547829e-11, 
    2.185843e-10, -1.289045e-10, 7.712231e-11, 1.131426e-09, -5.808531e-09, 
    7.884324e-10, 2.425651e-10, 7.423751e-11, 4.732148e-11, 5.115552e-10, 
    -8.093082e-10, -5.903217e-10, -3.706901e-11, -1.784173e-11, 9.443539e-10, 
    -2.337543e-10, -3.021143e-10, 8.915606e-10, 1.024034e-10, -4.828848e-12, 
    -9.056151e-10, 9.763248e-10, -4.655298e-11, 1.697096e-10, -2.215273e-09, 
    -2.826042e-09, -3.071563e-09, -3.507481e-09, -1.068884e-09, 4.311502e-09, 
    7.88873e-10, -4.227161e-10, 2.441851e-10, -1.677449e-10, -8.603251e-11, 
    3.020944e-11, 1.173497e-10, 6.79945e-12, -4.697931e-11, -8.078871e-11,
  -1.340315e-09, -1.909687e-09, 2.158711e-09, -1.758398e-09, 9.192114e-10, 
    -1.853263e-08, 3.240185e-09, -1.049077e-09, 2.238718e-09, 3.899398e-09, 
    2.771937e-09, 5.040445e-09, 2.01819e-10, -3.584013e-10, -8.801102e-10, 
    1.706943e-10, -2.072833e-09, 3.008118e-10, 1.319833e-11, 4.949605e-10, 
    -1.106777e-10, -2.618812e-10, -1.762501e-11, 1.825665e-09, -3.93047e-09, 
    -3.610925e-09, 9.744209e-09, -1.384206e-08, 4.871392e-09, 2.498211e-08, 
    -8.356441e-09, -4.554384e-09, 3.109985e-09, 1.666049e-09, 2.776765e-10, 
    -2.881652e-09, 3.101938e-10, 3.525358e-11, -7.280992e-09, 1.171065e-09, 
    -2.878816e-09, -5.464678e-10, 1.302727e-09, -3.644733e-10, 3.747935e-10, 
    -4.506582e-10, 1.901093e-10, 1.832145e-09, -1.249115e-09, -9.789325e-11, 
    5.907879e-10, -1.412165e-09, -1.46107e-09, 4.321087e-10, 1.047538e-09, 
    6.36291e-12, -1.986997e-10, 9.213607e-12, 3.050777e-09, -1.16173e-09, 
    -7.077361e-11, -2.841638e-10, 1.080558e-10, 6.343861e-10, -9.513804e-10, 
    1.122094e-08, -1.189168e-09, 3.915542e-09, -1.769966e-09, -3.265772e-09, 
    -3.429399e-10, 1.981737e-08, 4.763159e-10, -1.796938e-09, -4.37948e-10, 
    1.966427e-11, 8.743228e-12, 1.324576e-09, 4.838512e-11, -1.420464e-09, 
    4.666099e-10, 5.848688e-11, 1.525784e-10, 3.452495e-09, 4.285024e-09, 
    -4.61629e-10, 1.496286e-09, 8.702372e-11, 4.167244e-10, 8.126726e-10, 
    -1.192266e-09, -4.978326e-10, -6.125234e-11, -1.45835e-09, -1.899174e-10, 
    -2.252229e-10, -3.071968e-10, 1.701462e-09, 8.16236e-11, 6.052332e-11, 
    4.7336e-10, 2.450019e-09, -6.90985e-11, 1.749321e-10, -3.620617e-09, 
    -1.157961e-09, -2.267175e-09, -4.562114e-09, -1.048821e-09, 5.926889e-09, 
    1.527692e-09, -4.800178e-10, 6.935998e-10, -8.878409e-10, -2.350511e-10, 
    4.481464e-11, 2.187548e-10, 3.188294e-11, -1.211777e-10, -9.612577e-11,
  -4.426965e-10, 2.974872e-09, -1.998671e-09, -1.6949e-09, -5.840121e-09, 
    -1.349741e-08, -4.983605e-09, -1.845194e-09, 1.761578e-09, 5.54769e-09, 
    3.185363e-09, 4.789882e-09, 1.470255e-10, -1.443226e-09, -1.108504e-09, 
    -8.132359e-10, -3.864252e-09, 4.020109e-10, -9.12479e-11, 1.039695e-09, 
    6.849632e-11, -3.444995e-10, -2.009415e-10, 2.282519e-09, -4.112962e-09, 
    2.860077e-10, 8.954828e-09, -1.248614e-08, 6.218755e-09, 5.153441e-08, 
    -1.236606e-08, -7.640409e-09, 8.588472e-10, 2.710948e-09, 4.912977e-10, 
    -7.781779e-09, 4.439471e-11, 5.776002e-11, -1.789661e-08, 1.547605e-09, 
    -5.229646e-09, -9.931682e-10, 1.386553e-09, -3.286913e-10, -5.685479e-10, 
    -3.231833e-10, 3.005169e-10, 3.20415e-09, -1.518703e-09, -1.868887e-10, 
    7.368008e-10, -1.904993e-09, -2.860699e-09, 5.223796e-10, 1.939203e-09, 
    -2.279421e-11, -1.835303e-09, -1.293188e-12, 3.226492e-09, -1.63673e-08, 
    3.274181e-10, -4.790763e-10, 4.997105e-10, -7.228778e-10, -5.518774e-09, 
    1.792978e-08, -3.244111e-09, 3.019096e-09, -9.225118e-10, -4.943274e-09, 
    -4.215792e-10, 1.73867e-08, 4.507683e-10, -9.085568e-10, -4.0824e-09, 
    -1.560352e-11, -4.959588e-11, 1.728942e-09, 4.763265e-11, -3.114565e-09, 
    6.545946e-10, 1.943157e-10, 1.868159e-10, 7.84334e-09, 7.979821e-09, 
    -6.378116e-10, 2.948155e-09, 1.146816e-10, 7.111294e-10, 1.251593e-09, 
    -5.023537e-10, -1.032186e-09, -1.038813e-10, -8.230281e-09, 
    -3.314824e-10, -7.300401e-11, -5.680363e-11, 9.189023e-10, 5.38023e-11, 
    1.93603e-10, 1.466873e-09, 3.932081e-09, -9.107737e-11, 1.124665e-10, 
    -1.804324e-09, 1.899991e-10, -2.391062e-09, -4.256037e-09, -1.763453e-09, 
    6.230863e-09, 1.936513e-09, -3.879563e-10, 1.434643e-09, -2.560142e-09, 
    -4.652634e-10, -7.162271e-13, 3.553424e-10, 7.243095e-11, -1.595541e-10, 
    -2.027889e-10,
  2.087518e-09, 3.355296e-09, 1.09651e-09, 6.891128e-10, -3.857934e-09, 
    -3.633801e-09, -1.876779e-08, 1.425434e-09, 4.925482e-10, 4.550969e-09, 
    4.182851e-09, 5.638441e-09, 1.422222e-10, 5.940137e-10, -6.088214e-10, 
    -3.691896e-10, -2.491962e-09, -9.241319e-10, 2.043841e-10, 1.946233e-09, 
    1.98952e-13, -4.802985e-10, -2.766569e-10, 9.573853e-10, 3.217792e-09, 
    6.453035e-09, 2.294684e-08, -1.732926e-08, 1.0766e-08, 3.12312e-08, 
    -1.591658e-08, -6.209177e-09, -1.442771e-09, 3.491039e-09, 2.815739e-10, 
    -1.057163e-08, -5.101725e-10, 5.539391e-11, -1.604892e-08, 2.301132e-09, 
    -7.220575e-09, -1.566747e-09, 1.638519e-09, -6.223124e-10, -7.071321e-11, 
    -7.991616e-10, 2.993374e-10, 4.614748e-09, -9.217274e-10, -2.523404e-10, 
    1.520959e-09, -1.645191e-09, -4.783115e-09, 6.167681e-10, 2.927072e-09, 
    -8.442669e-11, -3.964345e-09, 4.16776e-11, 1.22412e-09, -2.677485e-08, 
    1.834479e-09, -6.336904e-10, 3.628315e-10, -3.940937e-09, -8.918613e-09, 
    2.193494e-08, -2.639638e-09, 2.055515e-09, -4.139991e-09, -6.123969e-09, 
    3.307719e-10, 1.334342e-09, 1.541594e-10, 2.008107e-09, -5.306108e-09, 
    -6.335199e-11, -1.361613e-10, 2.021743e-09, 2.017444e-11, 4.068056e-09, 
    -2.607123e-10, 2.774305e-10, 1.800089e-10, 7.160594e-09, 6.524033e-09, 
    5.994139e-11, 2.317165e-09, 1.712408e-10, 1.433352e-09, 2.354042e-09, 
    2.968875e-09, -3.383894e-09, -2.014318e-10, -2.016088e-08, 1.117883e-09, 
    1.71201e-10, 2.34121e-10, -1.798867e-09, -7.941026e-11, 1.487763e-10, 
    2.917943e-09, 4.658505e-09, -7.474021e-11, 4.03908e-11, -1.724061e-10, 
    3.343246e-10, -1.218723e-10, 9.634959e-11, -3.353165e-09, 3.86575e-09, 
    1.123055e-09, 1.073488e-10, 2.452822e-09, -3.613167e-09, -5.085496e-10, 
    -6.776872e-11, 3.55687e-10, 1.225953e-10, -1.521627e-10, -3.431637e-10,
  5.588561e-09, -2.569095e-09, 1.918465e-10, 1.543867e-09, 2.204843e-09, 
    2.007255e-09, -1.501502e-08, 3.954312e-09, 4.86466e-10, 2.567162e-09, 
    2.506169e-09, 4.228468e-09, 1.651756e-09, 1.511751e-09, 3.373088e-09, 
    -2.072244e-09, -2.785708e-09, -2.188301e-09, -1.849969e-10, 2.5438e-09, 
    -8.87951e-10, -2.368665e-10, -2.851834e-10, 1.79341e-10, 2.779984e-09, 
    7.378958e-09, 2.976401e-08, -3.325857e-08, 1.936513e-08, -1.9254e-09, 
    -2.14788e-08, -4.337267e-09, -4.633421e-09, 4.318451e-09, 4.444018e-10, 
    -1.211367e-08, -1.255637e-09, 6.012613e-11, 2.543175e-09, 3.884896e-09, 
    -1.098144e-08, -2.697789e-09, 2.424926e-09, -1.30981e-09, 5.141032e-09, 
    -6.574908e-09, 5.31287e-10, 6.272089e-09, 7.611675e-10, -4.316085e-10, 
    3.318874e-09, -1.272724e-09, -8.223997e-09, 5.31361e-10, 3.262612e-09, 
    -1.046772e-10, 1.924718e-10, 2.134755e-10, -1.512251e-09, -1.896744e-08, 
    6.101175e-09, -2.589218e-10, -1.304272e-09, -1.412138e-09, -5.244533e-09, 
    2.732384e-08, -2.2672e-09, 3.851994e-09, -2.719844e-09, -6.483958e-09, 
    1.728665e-09, 1.463383e-08, -1.729006e-09, -4.570779e-10, -4.340501e-09, 
    -1.817284e-10, -2.488676e-10, 2.716817e-09, -5.028511e-11, 1.558095e-08, 
    -2.826255e-10, 6.647136e-10, 2.194156e-10, 4.749722e-09, 2.603997e-09, 
    3.63957e-09, 2.750653e-10, 2.805791e-10, 2.345533e-09, 4.062628e-09, 
    7.790049e-09, -6.215089e-09, -2.695657e-10, -2.836356e-08, -4.371259e-10, 
    5.47584e-10, -1.597493e-09, -4.806793e-09, -2.00771e-10, -9.238193e-11, 
    1.798185e-09, 5.857824e-09, -1.005169e-10, -1.673328e-12, -7.622134e-10, 
    4.932303e-10, 8.81812e-10, 2.499462e-09, -2.564207e-10, 4.318053e-09, 
    1.418869e-09, 4.226877e-10, 2.840977e-09, -4.239553e-09, -3.011564e-10, 
    -1.056662e-10, 3.328324e-10, 1.065565e-10, -1.341078e-10, -5.832135e-10,
  9.005248e-09, -3.317211e-09, 1.26073e-09, -6.505729e-10, 4.53042e-11, 
    3.415153e-10, -1.235037e-09, 1.598892e-09, 9.989094e-10, 8.221832e-10, 
    1.346507e-09, 3.56016e-09, 2.663171e-09, -3.430046e-09, 8.085522e-09, 
    8.904864e-10, -6.779942e-10, -3.421889e-09, -1.537153e-09, 2.356785e-09, 
    3.045386e-09, 6.573373e-10, -1.814442e-10, 7.12248e-11, -1.452349e-09, 
    4.287472e-09, 1.827294e-08, -6.253532e-08, 3.106999e-08, -9.928783e-09, 
    -2.533108e-08, -3.44744e-09, -4.420087e-09, 5.448044e-09, 1.95206e-09, 
    -2.08255e-08, -1.440338e-09, 5.059064e-12, 1.259872e-08, 6.599987e-09, 
    -2.07991e-08, -4.788205e-09, 3.054311e-09, -2.658883e-09, 9.771668e-09, 
    -9.936457e-09, 1.040206e-09, 8.39357e-09, 3.041464e-09, -4.107257e-10, 
    6.691145e-09, 2.711431e-11, -1.335435e-08, 3.766559e-10, 2.593413e-09, 
    -3.052492e-11, 4.302535e-09, 4.208801e-10, -4.418979e-09, -4.147068e-09, 
    1.510159e-08, 9.433165e-10, -2.520324e-09, 6.087202e-09, -9.780808e-09, 
    1.572602e-08, -2.005891e-09, 6.750724e-09, 2.415106e-09, -4.606079e-09, 
    1.7194e-09, 4.249438e-08, -2.574325e-09, 1.953708e-10, 2.70129e-09, 
    -3.169589e-10, -3.401652e-10, 4.269467e-09, -1.11568e-10, 2.214358e-08, 
    6.847074e-10, 1.588349e-09, 4.075957e-10, -3.716252e-09, 7.476615e-10, 
    4.23961e-09, -3.813625e-09, 2.832508e-10, 3.293197e-09, 5.951648e-09, 
    9.746941e-09, -8.285542e-09, -8.870416e-11, -1.622169e-08, 5.470611e-10, 
    9.694304e-10, -7.859615e-09, -1.194456e-08, -7.787548e-11, -5.133871e-10, 
    -1.834906e-10, 6.962427e-09, -2.34408e-10, -6.412293e-11, -5.302127e-09, 
    5.204583e-10, 6.742766e-10, 7.475478e-10, -1.080707e-09, 1.127751e-08, 
    5.048093e-09, 4.721414e-10, 2.625768e-09, -5.450431e-09, -1.504645e-09, 
    -8.922143e-11, 1.65592e-10, 4.961365e-11, -1.169127e-10, -5.067591e-10,
  1.116376e-08, -1.009766e-09, 2.520324e-09, -6.23686e-10, -1.819899e-09, 
    -1.633737e-09, 3.219668e-09, -7.853544e-09, 9.223413e-10, 4.954472e-10, 
    -4.791332e-10, 1.204398e-09, 2.967397e-09, -1.195025e-08, 5.489312e-09, 
    9.687257e-11, -8.616325e-10, -3.524917e-09, -3.02304e-09, 1.793239e-09, 
    8.543338e-09, -8.48388e-10, 3.817604e-10, -5.836682e-10, -1.683247e-09, 
    -2.835463e-09, 7.861274e-09, -7.553183e-08, 1.835303e-08, -2.665331e-09, 
    -2.06345e-08, -3.99325e-09, -4.974424e-09, 7.554092e-09, 5.544621e-09, 
    -3.302677e-08, -1.799253e-09, -4.167333e-11, -1.557919e-08, 1.176958e-08, 
    -3.816076e-08, -5.228458e-09, 3.942688e-09, -4.461303e-09, 7.185008e-09, 
    -1.101512e-08, 1.903288e-09, 1.22572e-08, 5.637844e-09, -4.420784e-10, 
    9.661036e-09, 6.355094e-10, -2.176361e-08, -4.437198e-11, 2.291336e-09, 
    8.461143e-11, 9.047994e-09, 1.831552e-10, -8.693275e-09, 3.298375e-09, 
    2.177376e-08, 2.177785e-09, -3.572211e-09, 1.300888e-08, -1.313949e-08, 
    5.442701e-09, 1.155513e-09, 9.67492e-09, 2.702507e-09, 2.615934e-10, 
    9.437144e-10, 8.061841e-08, -5.758807e-10, 5.249944e-09, 1.645004e-08, 
    -5.119887e-10, -2.958842e-10, 6.992664e-09, -1.728324e-10, 2.748641e-08, 
    1.802363e-09, 2.520665e-09, 7.158292e-10, -3.390085e-09, 2.695685e-09, 
    2.516572e-09, -5.011088e-09, 1.980993e-10, 3.220753e-09, 8.161607e-09, 
    8.526456e-09, -6.914457e-09, 8.775487e-10, 1.00538e-08, 2.034199e-09, 
    1.355892e-09, -1.558374e-08, -2.421655e-08, 1.435865e-10, -9.904625e-10, 
    3.050786e-10, 4.760459e-09, -3.960601e-10, -3.031353e-10, -1.689409e-08, 
    -1.17484e-09, 1.392777e-09, -3.744674e-09, -2.174204e-09, 1.52466e-08, 
    5.657398e-09, -1.454737e-09, 2.583079e-09, -6.219523e-09, -5.942411e-09, 
    -5.114202e-11, -7.165113e-11, 8.025225e-11, -1.087805e-10, 5.798029e-12,
  9.090513e-09, -8.761845e-10, 1.569674e-09, 4.91525e-10, -1.189733e-09, 
    -2.33814e-09, -2.888896e-09, -1.891487e-08, -5.216521e-10, 2.484796e-09, 
    -1.417561e-09, 1.982698e-10, -1.348894e-09, -5.048491e-09, -7.187282e-09, 
    -2.141792e-09, -4.08815e-09, -2.029822e-09, -4.008591e-09, 1.630497e-09, 
    1.273781e-08, -2.290335e-09, 3.936407e-10, -4.198455e-10, 4.454819e-10, 
    -2.64879e-09, 1.808723e-08, -8.557367e-08, 2.037041e-09, -2.99957e-09, 
    -1.467617e-08, -6.167795e-09, -6.851792e-09, 8.428174e-09, 6.946948e-09, 
    -3.878262e-08, -2.739841e-09, -1.201528e-11, -6.115499e-08, 2.109548e-08, 
    -5.773502e-08, 1.757883e-09, 5.110522e-09, -6.616418e-09, -2.412776e-09, 
    -5.589015e-09, 1.948138e-09, 2.066966e-08, 8.003019e-09, -3.530367e-10, 
    1.109702e-08, -1.239073e-09, -3.282078e-08, -2.856951e-11, 3.496258e-09, 
    1.841158e-10, 1.103456e-08, -1.299782e-09, -7.002569e-09, 5.777864e-09, 
    8.448126e-09, 3.155321e-09, -1.719343e-09, 1.392565e-08, -9.129622e-10, 
    1.441651e-08, 6.105722e-09, 1.618412e-08, 7.874348e-09, -2.059323e-09, 
    -1.275964e-09, 3.48324e-08, 4.343406e-10, 2.701711e-09, 2.674655e-08, 
    -7.779022e-10, -2.236007e-10, 1.147927e-08, -4.243987e-10, 3.206435e-08, 
    1.15827e-09, 2.489863e-09, 1.18203e-09, -2.4786e-09, 4.38979e-09, 
    2.128786e-10, -1.578712e-09, -1.153921e-10, 1.742846e-09, 7.897597e-09, 
    8.224958e-09, -4.863432e-09, 2.069967e-09, 3.835934e-08, 2.616105e-09, 
    1.416157e-09, -1.874473e-08, -2.00954e-08, 4.860112e-10, -1.484545e-09, 
    1.877538e-10, 1.223086e-09, -1.036483e-09, -8.625491e-10, -2.323674e-08, 
    1.816886e-09, 5.779214e-09, -6.796597e-09, 7.322228e-09, 1.656457e-08, 
    3.930722e-09, -2.441709e-09, 2.245372e-09, -6.912444e-09, -7.343999e-09, 
    -2.677325e-12, -3.511929e-10, 2.869882e-11, -1.01938e-10, 1.22435e-09,
  5.409447e-09, -1.456783e-09, -5.344987e-10, -1.419266e-09, -1.274657e-09, 
    -3.438856e-09, -1.006708e-08, -1.534897e-08, -3.297373e-09, 1.543697e-09, 
    1.103842e-09, -2.203876e-09, -3.912191e-09, 8.701647e-09, -8.322274e-09, 
    -4.510849e-09, -6.743557e-09, 9.519283e-10, -5.696009e-09, 2.463082e-09, 
    1.721179e-08, 7.028859e-09, -2.757247e-09, 4.831691e-10, 1.970591e-09, 
    -6.071446e-10, -6.85373e-08, -6.125521e-08, -2.409394e-08, -3.633318e-09, 
    -2.206042e-08, -8.254688e-09, -7.910387e-09, 7.49759e-09, 4.039123e-09, 
    -5.849472e-08, -3.806627e-09, 6.712497e-11, -7.600181e-08, 3.750071e-08, 
    -7.708888e-08, 9.261385e-09, 5.940052e-09, -1.086532e-08, -2.267899e-08, 
    1.08389e-08, -3.535519e-09, 3.205137e-08, 1.004937e-08, -2.831051e-10, 
    1.005132e-08, -7.83848e-09, -4.948288e-08, 6.124307e-11, 4.540128e-09, 
    2.550564e-10, 7.859796e-09, -4.632363e-09, 3.245719e-09, -7.697416e-09, 
    -1.192757e-08, 2.782372e-09, -8.230927e-11, 1.178946e-08, 2.691683e-09, 
    2.01897e-08, 1.982988e-08, 6.303083e-08, 1.473546e-08, -4.368587e-09, 
    -5.617153e-09, -1.195133e-08, -1.250015e-08, -7.692051e-10, 2.531248e-08, 
    -1.059789e-09, -1.386056e-10, 1.598707e-08, -8.851572e-10, 2.715484e-08, 
    -2.989054e-09, 9.599042e-10, 1.838345e-09, 2.960974e-10, 1.83644e-09, 
    -1.147328e-09, -5.516654e-10, -1.117655e-09, -1.727258e-10, 6.827605e-09, 
    8.777477e-09, -2.781769e-09, 3.020062e-09, 3.909047e-08, 7.820518e-10, 
    9.306462e-10, -1.699885e-08, 7.691767e-09, 2.514184e-10, -1.919159e-09, 
    6.477876e-10, 1.24448e-10, -1.885727e-09, -1.735089e-09, 9.047028e-09, 
    3.769117e-09, 2.934485e-09, -1.270962e-09, 1.438542e-08, 1.058538e-08, 
    1.512205e-09, -4.542073e-09, -6.700702e-10, -8.155496e-09, -6.124083e-09, 
    6.263007e-11, 3.811351e-10, 2.037126e-11, -6.379608e-11, 4.38456e-09,
  1.558135e-09, -1.294893e-10, 7.593144e-10, -3.092453e-09, -1.106457e-09, 
    -2.921411e-09, -1.096009e-08, -1.737192e-09, -1.279034e-08, 
    -2.996728e-09, 5.356924e-10, -2.822105e-09, 1.906983e-09, 1.080855e-08, 
    9.113251e-09, -6.857237e-09, -8.495317e-09, 4.261835e-09, -7.659892e-09, 
    3.712216e-09, 1.690267e-08, 5.772904e-09, -1.069168e-09, 7.632366e-10, 
    2.772367e-09, 6.8394e-10, -5.557609e-08, -2.395001e-08, -4.997679e-08, 
    1.252403e-08, -2.225676e-08, -1.102887e-08, -6.228277e-09, 5.322534e-09, 
    4.7919e-10, -6.785683e-08, -4.269759e-09, 1.237268e-10, -6.414012e-08, 
    6.271726e-08, -8.737933e-08, 6.754419e-09, 6.690826e-09, -1.813859e-08, 
    8.282655e-10, 2.545238e-08, -1.005418e-08, 4.699395e-08, 1.21909e-08, 
    -3.607354e-10, 7.641212e-09, -1.582345e-08, -6.805185e-08, -3.029982e-10, 
    4.565211e-09, 2.714273e-10, -3.657249e-09, -6.705056e-09, 1.754191e-08, 
    -1.579234e-08, -3.012246e-09, 6.832011e-10, -1.780336e-10, 1.278996e-08, 
    -3.180446e-09, 2.340124e-08, 3.670596e-08, 5.100406e-08, 1.808337e-08, 
    -2.627644e-09, -4.094522e-08, -4.741065e-08, -5.161098e-09, 
    -2.653735e-09, 1.46007e-08, -1.233161e-09, 2.994724e-10, 1.867403e-08, 
    -1.820115e-09, 1.582356e-08, 3.05505e-10, -5.785097e-10, 2.827392e-09, 
    7.286189e-10, 1.090257e-10, -2.016066e-09, -3.254286e-09, -1.723549e-09, 
    -1.181167e-09, 7.499665e-09, 4.337267e-09, 6.264076e-09, 3.729852e-09, 
    -8.570578e-09, -1.442686e-09, -3.581133e-13, -1.732089e-08, 7.558867e-09, 
    -2.050172e-09, -2.077672e-09, 2.887646e-10, -8.678285e-10, -2.556558e-09, 
    -2.826084e-09, 6.486005e-09, 1.324509e-09, -3.069545e-12, 2.757247e-09, 
    8.480697e-09, 2.711658e-09, -3.431467e-09, -4.17765e-09, -1.635044e-09, 
    -9.767746e-09, -1.235793e-08, 1.519879e-10, 9.375469e-10, 2.903278e-11, 
    -3.523937e-11, 5.956792e-09,
  2.781917e-10, -2.847855e-11, 3.696925e-09, -1.250555e-10, -1.478725e-09, 
    -1.025342e-09, -8.380368e-09, 1.076654e-08, -2.582368e-08, -1.029974e-08, 
    -4.042136e-09, -6.02995e-10, 2.864738e-09, 4.301171e-09, 1.908643e-08, 
    -1.835798e-09, -9.984598e-09, 8.267762e-09, -1.171262e-08, 3.07034e-09, 
    1.290647e-08, -2.870593e-11, 1.923809e-09, -1.347473e-09, 3.099501e-09, 
    1.346621e-09, 2.662688e-08, -1.800936e-08, -1.126881e-07, 2.913316e-08, 
    -2.524536e-08, -9.387293e-09, -4.871879e-09, 2.783395e-09, 2.47195e-09, 
    -7.25193e-08, -2.078548e-09, 4.206768e-10, -4.763143e-08, 9.055879e-08, 
    -9.453464e-08, 3.39827e-09, 7.374851e-09, -2.722733e-08, 1.26488e-09, 
    1.811037e-08, -1.010989e-08, 6.58127e-08, 1.506426e-08, -5.499068e-10, 
    -1.937693e-09, -1.048397e-08, -8.355227e-08, -5.033712e-10, 5.141662e-09, 
    1.084857e-10, -3.380001e-08, -1.486852e-08, 2.668394e-08, -6.892904e-10, 
    1.278414e-08, 1.208377e-09, -1.304954e-09, 1.472475e-08, -9.177962e-09, 
    3.171698e-08, 1.249905e-07, 8.857853e-09, 1.352595e-08, -1.338265e-09, 
    -7.631581e-08, -6.392668e-08, 9.254109e-10, -4.054755e-09, 8.670634e-09, 
    -9.493419e-10, 1.515446e-10, 1.95564e-08, -3.077054e-09, 5.276377e-09, 
    -3.315876e-09, 1.723279e-09, 4.317684e-09, 1.191154e-09, -1.858211e-09, 
    -2.335696e-09, -3.336993e-09, 1.732019e-10, -3.966392e-10, 1.340302e-08, 
    7.848371e-10, 1.95973e-08, 3.398398e-09, -1.198072e-07, -9.371774e-10, 
    -1.124806e-09, -2.599634e-08, 2.099125e-08, -5.660979e-09, -2.089632e-09, 
    -4.909566e-10, 1.81862e-09, -2.794255e-09, -3.716416e-09, -2.433524e-09, 
    -1.821775e-09, 3.591936e-09, 2.889351e-09, 2.550905e-09, -6.536993e-11, 
    -5.90893e-09, -1.315357e-09, -9.243877e-10, -9.73489e-09, -1.421193e-08, 
    2.365709e-10, 1.260531e-09, 5.823075e-11, 3.801404e-13, 7.103552e-09,
  -2.420279e-09, -4.984599e-10, -2.398963e-09, 2.1924e-08, -5.741185e-10, 
    8.50946e-10, -4.454705e-09, 9.848918e-09, -2.977839e-08, -1.431101e-08, 
    -4.660308e-09, 4.359549e-09, 8.506618e-10, 2.767763e-09, 3.783663e-08, 
    7.986285e-09, -1.446597e-08, 1.176809e-08, -1.45971e-08, -7.712515e-10, 
    1.247298e-08, 1.170633e-09, 1.292563e-09, -6.25846e-10, 2.170623e-09, 
    -8.628831e-11, 6.192408e-09, -1.673334e-08, -9.803773e-08, 2.744298e-08, 
    -2.880699e-08, -2.757929e-09, -5.341008e-09, 8.903669e-09, 1.333024e-08, 
    -7.89222e-08, 1.178006e-09, 1.000288e-09, -2.599751e-08, 1.154747e-07, 
    -7.904411e-08, 4.023889e-09, 7.057551e-09, -3.456545e-08, -1.583311e-08, 
    1.26077e-08, -5.977e-09, 9.04588e-08, 1.859178e-08, -7.684378e-10, 
    -9.709119e-09, -8.65623e-09, -1.017782e-07, -1.240778e-09, 7.96121e-09, 
    -1.300862e-10, -7.662283e-08, -2.825556e-08, 1.639521e-08, 2.768206e-08, 
    8.792995e-09, 1.929209e-09, -2.549996e-10, 1.689807e-08, -1.033989e-08, 
    3.999531e-08, 1.364933e-07, 6.305402e-08, 9.197095e-09, -3.887408e-09, 
    -8.256495e-08, -3.279354e-08, 3.587218e-09, -2.887987e-09, 1.671915e-08, 
    -1.097646e-10, 9.136158e-11, 1.734414e-08, -4.646729e-09, -1.850822e-10, 
    -5.936073e-09, 9.963557e-09, 6.21452e-09, 1.278977e-11, -4.012122e-09, 
    -2.611841e-09, 3.314369e-09, 4.957656e-09, -1.309754e-09, 1.29653e-08, 
    -5.156835e-10, 2.668121e-08, 2.325038e-09, -1.603801e-07, -6.971277e-09, 
    -1.749493e-09, -3.728361e-08, 4.965278e-08, -8.773384e-09, -2.976754e-09, 
    2.837623e-10, 2.275531e-09, -2.551769e-09, -3.471918e-09, -4.128765e-09, 
    -3.378489e-09, 7.350593e-09, 9.81305e-09, 1.790511e-09, -1.350827e-09, 
    -5.915183e-09, 1.206104e-09, -1.324395e-09, -8.355244e-09, -2.252364e-09, 
    2.098204e-10, 1.849848e-09, 1.468337e-10, 7.000622e-11, 7.716949e-09,
  -5.976801e-09, 4.12399e-10, -6.880725e-09, 5.552403e-08, 4.918661e-10, 
    6.322693e-10, -2.160789e-09, -2.586887e-09, -1.402003e-08, -9.703797e-09, 
    -9.723067e-10, 6.254652e-09, -5.742891e-10, 1.127205e-10, 2.051087e-08, 
    -7.655956e-09, -1.634623e-08, 1.550461e-08, -1.891695e-08, -5.039567e-09, 
    1.248492e-08, -2.523336e-09, -5.470042e-10, 5.191339e-09, -5.188099e-10, 
    -1.847923e-09, -3.081425e-09, -1.466566e-08, -3.97377e-08, 1.866169e-10, 
    -3.900237e-08, 1.303334e-08, 7.436648e-08, 1.468078e-08, 2.630571e-08, 
    -8.075125e-08, 4.287392e-09, 2.038107e-09, -1.172964e-09, 1.316288e-07, 
    -6.950835e-08, 4.82413e-09, 9.464003e-09, -3.348412e-08, -5.467484e-09, 
    -5.038163e-08, -6.844402e-09, 1.246964e-07, 1.845616e-08, -1.253795e-09, 
    -1.421851e-08, -5.591886e-08, -1.094346e-07, 2.319177e-09, 1.349575e-08, 
    -5.018705e-10, -1.144388e-07, -3.653248e-08, -2.696631e-08, 5.287349e-08, 
    -3.916682e-09, 7.633503e-10, 1.470596e-09, 1.623502e-08, -2.255422e-09, 
    5.77748e-08, 1.11294e-07, 3.705389e-08, 1.758048e-08, -4.265132e-09, 
    -7.655018e-08, 2.384525e-09, -2.385281e-08, 1.847354e-09, 2.332134e-08, 
    1.264596e-09, 9.852101e-10, 1.509838e-08, -6.104995e-09, -7.174208e-10, 
    -8.181132e-09, 2.538027e-08, 7.680342e-09, -2.243326e-09, 5.59055e-10, 
    2.718991e-09, 9.470966e-09, 6.506355e-09, 5.410875e-09, -2.793286e-10, 
    -1.126352e-09, 2.235857e-08, 4.502567e-10, -1.489845e-07, -1.757525e-08, 
    -1.904016e-09, -4.811258e-08, 5.633177e-08, -1.26285e-08, -6.004041e-09, 
    1.757996e-09, 4.801706e-10, -2.605653e-09, -1.998757e-09, -4.221135e-09, 
    -6.476569e-09, 6.782045e-09, 1.727966e-08, 4.55799e-09, -1.200704e-09, 
    -4.828564e-09, 1.660339e-09, -1.216961e-09, -5.449408e-09, 5.137565e-09, 
    1.181888e-10, 2.502304e-09, 1.950227e-10, 1.451781e-10, 6.179619e-09,
  -6.269545e-09, 2.168406e-09, 3.979039e-13, 8.887883e-08, 1.721276e-09, 
    -1.695241e-09, -2.080299e-09, -4.538322e-09, 1.099028e-08, 5.172183e-10, 
    7.892538e-09, 3.736034e-09, -4.028493e-10, -1.369187e-09, -5.160814e-10, 
    -6.259582e-08, -1.217322e-08, 2.174306e-08, -3.054537e-08, -2.800732e-09, 
    7.783854e-09, -8.253096e-10, -2.271389e-08, -6.396988e-09, -6.33969e-09, 
    -6.357311e-09, -9.383513e-08, -1.28943e-08, -3.00401e-08, -1.363031e-08, 
    -7.418527e-08, 1.377185e-08, -1.693417e-08, 1.221457e-08, 4.45844e-08, 
    -7.508032e-08, 7.526785e-09, 2.720114e-09, 2.840437e-08, 1.340845e-07, 
    -6.251584e-08, 4.890978e-09, 1.631892e-08, -2.476056e-08, -5.678146e-09, 
    -1.149168e-07, -1.074307e-08, 1.663334e-07, 9.154462e-09, -1.803407e-09, 
    -1.560508e-08, -1.119897e-07, -1.084623e-07, 6.62493e-09, 1.981808e-08, 
    -6.456276e-10, -1.416097e-07, -4.097527e-08, -1.054298e-07, 6.241584e-08, 
    -9.057999e-10, 7.47491e-11, 3.09393e-09, 1.039017e-08, 1.196291e-08, 
    6.40502e-08, 8.686521e-08, -5.515386e-08, 2.068765e-08, -4.162246e-09, 
    3.14742e-10, -3.379847e-08, -5.409032e-08, 2.265836e-09, 2.114568e-08, 
    3.082448e-09, 1.002263e-09, 8.421978e-09, -7.405566e-09, -2.776801e-10, 
    -5.69247e-09, 4.133176e-08, 8.142081e-09, -2.587001e-09, 9.525991e-09, 
    9.868302e-09, 1.305824e-08, 5.929849e-09, 3.198189e-08, -1.059709e-08, 
    -1.600313e-09, -3.036905e-09, -1.65673e-09, -1.667935e-07, -2.389896e-08, 
    1.361172e-10, -6.085017e-08, -2.889436e-08, -1.546329e-08, -1.056068e-08, 
    3.46688e-10, -6.861001e-11, -5.572907e-09, -3.65219e-12, 4.627225e-09, 
    -2.465043e-08, 1.902606e-09, 1.551683e-08, 1.025472e-08, -7.968879e-10, 
    -3.657817e-09, 8.603251e-10, -2.726779e-10, -1.073374e-09, 2.87713e-09, 
    1.942908e-11, 3.059569e-09, 2.520508e-10, 2.068319e-10, 3.831872e-09,
  -3.455159e-08, 1.17268e-09, 2.728484e-12, 1.299788e-07, -1.072067e-10, 
    -5.787228e-09, -8.290044e-10, -2.801471e-09, 1.939327e-08, 1.190756e-08, 
    1.09502e-08, 1.600938e-09, -4.905587e-10, -1.33507e-08, -2.584557e-09, 
    -1.28233e-07, -5.736537e-09, 2.872088e-08, -1.486885e-08, 1.170793e-08, 
    -2.43233e-09, -6.888285e-09, -1.110732e-08, -1.511296e-08, -1.255194e-08, 
    -3.81624e-09, -2.257455e-07, -1.600358e-08, -3.144771e-08, -6.697292e-09, 
    -1.158243e-07, -8.576455e-08, -3.411776e-08, 6.092705e-09, 6.954394e-08, 
    -6.910489e-08, 1.173347e-08, 3.306781e-09, 1.03455e-08, 1.272839e-07, 
    -6.6536e-08, 2.940965e-09, 1.909657e-08, -1.756195e-08, -2.995114e-08, 
    -5.508446e-08, 2.957847e-09, 2.08218e-07, -1.331596e-08, -2.39325e-09, 
    -1.241611e-08, -1.342927e-07, -1.112962e-07, 7.143512e-09, 2.303736e-08, 
    -7.552217e-10, -1.349529e-07, -7.498961e-08, -1.826721e-07, 6.849579e-08, 
    6.61862e-09, -5.707079e-11, 4.490403e-09, -2.328079e-09, 3.195671e-08, 
    7.497874e-09, 4.74231e-08, 1.868875e-08, 1.459318e-08, 7.005383e-10, 
    2.786271e-08, -9.644896e-08, -5.565744e-08, 5.416041e-10, 1.220088e-08, 
    3.12707e-09, 6.752572e-10, 5.574094e-09, -8.244496e-09, 7.85576e-10, 
    -3.478135e-09, 5.331783e-08, 8.931124e-09, -1.796252e-10, 1.089631e-08, 
    2.251909e-09, 1.265153e-08, 2.926527e-09, 6.481056e-08, -4.214826e-09, 
    -7.335075e-10, -6.374e-08, -1.840959e-09, -2.208889e-07, 1.841187e-07, 
    6.572691e-10, -7.301944e-08, 5.902052e-08, -1.926617e-08, -1.438113e-08, 
    -7.807216e-09, 3.325326e-09, -4.935295e-09, 1.861594e-09, 5.023674e-08, 
    -4.576168e-08, -2.019965e-08, 1.733792e-08, 2.046443e-08, -3.637069e-09, 
    -4.504727e-09, -5.725269e-10, 1.771241e-10, 1.935064e-09, 2.03886e-09, 
    -2.254069e-10, 3.458908e-09, -2.485478e-11, 2.296261e-10, 6.620439e-09,
  -3.27384e-08, 6.676828e-10, 1.820013e-09, 1.200078e-07, -2.247702e-09, 
    -1.09095e-08, 4.597496e-09, -6.646133e-09, 1.847104e-08, 4.43049e-09, 
    2.482579e-09, -6.662049e-10, -8.30255e-10, -7.256745e-08, -2.451543e-09, 
    -1.489759e-07, -6.377457e-09, 3.366546e-08, 3.629823e-08, 2.868001e-08, 
    -2.42751e-08, -7.446829e-09, -3.500759e-09, -1.299554e-09, 1.781814e-09, 
    4.977892e-09, -9.394864e-08, -2.321019e-08, -2.031504e-08, 4.174922e-09, 
    -1.327317e-07, -1.17631e-07, 9.239568e-08, -5.872141e-08, 6.433504e-08, 
    -7.428434e-08, 1.295713e-08, 3.27816e-09, -3.722448e-08, 1.07385e-07, 
    -6.021887e-08, 2.092634e-09, 1.504128e-08, -1.635342e-08, -6.674327e-09, 
    -1.809735e-08, 3.5065e-08, 2.383172e-07, -4.804883e-08, -5.036753e-09, 
    8.625548e-09, -9.973087e-08, -1.227472e-07, -2.441538e-10, 2.311012e-08, 
    -2.341892e-09, -1.090092e-07, -8.077825e-08, -1.751957e-07, 7.907926e-08, 
    4.876597e-09, -1.056151e-10, 1.410888e-08, -1.959679e-08, 5.214998e-08, 
    -3.341484e-08, 1.486092e-08, 3.446257e-08, 2.56797e-08, -6.729579e-09, 
    2.563115e-08, -1.32974e-07, -2.654428e-08, 3.086484e-09, 9.532733e-09, 
    -3.693003e-09, -5.025669e-10, -3.386361e-09, -8.159356e-09, 9.013888e-09, 
    -1.931596e-09, 5.986087e-08, 1.273264e-08, 1.159265e-09, -5.969923e-09, 
    8.054144e-09, -8.095981e-09, 5.110223e-10, 1.016049e-07, 6.66131e-09, 
    -3.575451e-10, -1.693833e-07, -1.693394e-09, -2.724635e-07, 1.886145e-07, 
    -4.887033e-09, -8.067775e-08, 5.365553e-08, -2.555817e-08, -1.746084e-08, 
    -5.447259e-08, 8.220582e-09, -2.604821e-09, 3.220961e-09, 7.150254e-08, 
    -6.937978e-08, -4.445133e-08, 1.349622e-08, 3.709658e-08, -2.478373e-11, 
    -5.998686e-09, -3.378659e-09, 1.694275e-09, 3.758487e-10, 4.52053e-09, 
    -4.156618e-10, 4.012975e-09, -2.749303e-10, 1.982343e-10, 2.162108e-08,
  -1.983324e-08, 7.836434e-10, 6.959908e-10, 5.393269e-08, -2.709442e-08, 
    -5.338507e-09, 1.224225e-08, -5.672518e-09, 1.022102e-08, 4.618983e-09, 
    -7.370318e-10, -3.638547e-09, 4.499725e-10, -1.182112e-07, -1.051012e-08, 
    -1.873931e-07, -3.629722e-09, 3.541362e-08, 2.17991e-08, 3.39171e-08, 
    -3.80611e-08, -1.362969e-08, 3.585683e-10, -4.18197e-09, 1.012086e-08, 
    4.936737e-09, -2.504146e-08, -1.795024e-08, -2.330819e-08, 1.044316e-08, 
    -1.163497e-07, -8.94579e-09, 1.409319e-08, -1.16561e-07, -6.148639e-09, 
    -8.764789e-08, 1.469688e-08, 3.47481e-09, -8.431346e-08, 8.347501e-08, 
    -4.536917e-08, 5.478341e-09, 1.684754e-08, -2.613099e-08, -5.11875e-09, 
    -4.043056e-08, 7.599897e-08, 2.384161e-07, -9.137311e-08, -8.736563e-09, 
    2.726397e-08, -8.533357e-08, -1.486961e-07, -3.401601e-09, 1.911993e-08, 
    -3.748255e-09, -1.06128e-07, -7.930065e-08, -1.018416e-07, 1.011343e-07, 
    -1.281478e-09, -1.286935e-10, 3.981779e-08, -3.568116e-08, 6.90701e-08, 
    -6.232688e-08, -9.078235e-09, 2.705804e-08, 3.113541e-08, -9.903033e-09, 
    2.122988e-09, -1.670072e-07, 6.967866e-09, -6.23686e-10, 9.918267e-09, 
    -1.042395e-08, -1.599631e-09, -5.973902e-09, -6.922974e-09, 2.549473e-08, 
    8.446023e-09, 5.426291e-08, 1.96776e-08, -1.036597e-09, -1.35484e-08, 
    1.584897e-08, 5.919288e-07, 4.798608e-09, 1.432234e-07, 4.477408e-08, 
    -2.244974e-09, -2.477452e-07, -2.502844e-09, -3.190906e-07, 2.409809e-08, 
    5.125275e-09, -7.978353e-08, 1.323565e-08, -2.787533e-08, -2.132242e-08, 
    -8.875963e-08, 3.194913e-09, 1.430504e-08, 3.444654e-09, 4.061212e-08, 
    -8.494328e-08, -3.608852e-08, 6.544497e-09, 5.723155e-08, 6.482878e-09, 
    -3.087621e-09, -6.799951e-09, 2.29204e-09, -2.736783e-09, 3.280093e-09, 
    -8.525831e-10, 4.397762e-09, -3.043752e-10, 1.350884e-10, 4.094932e-08,
  -3.491323e-10, 4.400817e-10, -5.828838e-09, 5.485617e-09, -3.186119e-08, 
    7.932613e-09, 1.728097e-08, 3.195623e-09, -6.016649e-09, -3.562945e-09, 
    -1.061949e-09, -1.498847e-09, 4.004164e-09, -3.598097e-08, -2.442096e-08, 
    -1.821757e-07, 1.399906e-08, 2.814204e-08, -3.404608e-09, 1.403328e-08, 
    -1.931801e-08, -2.198988e-08, 1.43848e-09, -1.766239e-09, 6.113851e-09, 
    -7.10088e-10, -3.131026e-08, -2.65527e-09, -4.699314e-08, 1.566798e-08, 
    -8.276049e-08, 3.582534e-08, -2.339561e-09, -9.407245e-09, -6.160587e-08, 
    -1.029661e-07, 1.781725e-08, 3.865864e-09, -1.044571e-07, 6.117872e-08, 
    -4.507131e-08, 1.052172e-08, 2.674187e-08, -3.00017e-08, -6.746404e-09, 
    -5.906327e-08, 9.076922e-08, 1.987638e-07, -1.252213e-07, -1.212789e-08, 
    3.677478e-08, -8.020049e-08, -1.766374e-07, -6.664322e-10, 1.330439e-08, 
    -4.454819e-10, -1.16932e-07, -7.936484e-08, -2.079723e-08, 1.19089e-07, 
    -3.778609e-09, -2.27044e-09, 5.541642e-08, -4.685232e-08, 8.022089e-08, 
    -5.717686e-08, -4.171886e-08, 2.744537e-08, 1.25508e-08, -1.487922e-08, 
    -2.747868e-08, -1.791002e-07, 4.011667e-08, 3.745868e-09, 1.507827e-08, 
    -4.146955e-09, -2.156497e-09, -1.304267e-08, -5.625574e-09, 4.112735e-08, 
    1.485398e-08, 3.42237e-08, 2.626143e-08, 1.230092e-09, -7.584049e-10, 
    2.090064e-08, 2.17146e-07, 1.763249e-08, 1.905098e-07, 1.403519e-07, 
    -1.431658e-09, -1.997466e-07, -2.848196e-09, -3.174414e-07, 
    -1.856188e-08, 1.362181e-08, -7.35014e-08, 8.416805e-09, -2.374156e-08, 
    -2.458489e-08, -8.083646e-08, -1.565991e-08, 4.272721e-09, 3.137124e-09, 
    4.380786e-08, -5.641607e-08, -1.683395e-08, -1.423666e-08, 7.565529e-08, 
    2.648085e-08, 5.380798e-10, -8.373263e-09, -1.650619e-09, -3.774062e-09, 
    -6.797336e-10, -1.202807e-09, 5.267935e-09, -4.671783e-10, 8.951417e-11, 
    4.285312e-08,
  5.587651e-09, 2.69722e-10, -5.666436e-09, -1.286907e-08, -1.214352e-08, 
    2.607743e-08, 2.141093e-08, 2.126916e-08, -9.517919e-09, -4.722722e-09, 
    -2.980698e-09, -2.767706e-10, 1.56337e-08, 1.215244e-07, -3.344593e-08, 
    -1.261799e-07, 1.700342e-08, -1.606571e-08, 2.706076e-08, -4.402324e-08, 
    2.437389e-09, -3.037047e-08, 2.757872e-09, -1.136243e-09, -7.998437e-10, 
    -4.336408e-08, -4.312312e-09, 1.467072e-09, -5.891565e-08, 2.675534e-08, 
    -6.650754e-08, 5.016824e-08, -1.022755e-08, 2.818848e-08, -4.339182e-08, 
    -1.030792e-07, 1.95176e-08, 2.923755e-09, -1.114349e-07, 4.210386e-08, 
    -2.185212e-08, 1.063262e-08, 1.802042e-08, -3.127293e-08, -2.257337e-08, 
    -6.328997e-08, 6.523368e-08, 1.336844e-07, -1.284865e-07, -1.519984e-08, 
    3.616147e-08, -7.051557e-08, -2.001166e-07, 5.378172e-09, 3.596242e-09, 
    -4.3201e-12, -1.301974e-07, -9.294136e-08, 4.008091e-08, 1.508732e-07, 
    1.68825e-11, -1.129939e-08, 3.704821e-08, -6.396557e-08, 7.151279e-08, 
    -4.082591e-08, -6.166528e-08, 2.583346e-08, -1.169218e-08, -2.311907e-08, 
    3.238628e-07, -1.139436e-07, 3.606959e-08, 1.191773e-08, 2.539282e-08, 
    4.843344e-09, -2.641869e-09, -2.065059e-08, -5.055046e-09, 2.461849e-08, 
    1.922518e-08, 1.656704e-08, 2.965322e-08, 3.296293e-09, 9.434132e-09, 
    2.983228e-08, -5.294163e-08, 2.929636e-08, 2.35367e-07, 2.012739e-07, 
    5.558661e-09, -1.047204e-07, -3.535462e-09, -3.199268e-07, -5.026703e-08, 
    -4.718425e-09, -4.346331e-08, 7.443526e-08, -9.518942e-09, -2.393168e-08, 
    3.247447e-08, -2.939182e-08, -1.611866e-09, 2.2942e-09, 6.057093e-08, 
    -5.001226e-08, -3.707277e-08, -1.677728e-08, 7.788066e-08, 4.435179e-08, 
    2.916636e-10, -8.978702e-09, -8.30056e-09, -3.217167e-09, -2.538229e-09, 
    -1.850242e-09, 6.666411e-09, -9.604442e-10, 9.576695e-11, -1.698578e-08,
  8.429254e-09, 1.262492e-10, -2.82688e-09, -9.775306e-09, -6.50806e-09, 
    3.676229e-08, 3.00742e-08, 6.133786e-08, -4.760466e-09, 9.566179e-10, 
    1.635328e-09, -2.475247e-09, 6.73964e-09, 5.517478e-08, 1.123965e-09, 
    -8.793718e-08, 1.342263e-08, 5.295442e-08, 7.860889e-08, -1.49611e-07, 
    2.451321e-08, -3.821282e-08, 3.029584e-09, -1.784315e-10, -2.040173e-08, 
    -1.090546e-07, -8.604445e-09, -5.444292e-09, -6.083172e-08, 1.196184e-08, 
    -8.78369e-08, 5.163128e-08, -1.72343e-08, 9.219377e-09, 9.538724e-09, 
    -8.37984e-08, 1.87918e-08, 2.420023e-09, -1.20656e-07, 2.213146e-08, 
    5.874574e-09, 1.170355e-08, -1.057504e-08, -3.518186e-08, -4.42131e-08, 
    -5.615146e-08, 1.285281e-08, 6.198076e-08, -1.07535e-07, -1.772336e-08, 
    3.274181e-08, -6.794272e-08, -2.118617e-07, 3.774141e-09, 1.504279e-09, 
    -4.296794e-10, -1.351144e-07, -6.920381e-08, 4.874436e-08, 2.114694e-07, 
    2.046875e-09, 1.359768e-08, 4.647603e-08, -7.42357e-08, 5.246581e-08, 
    -3.029908e-08, -5.231635e-08, 1.465008e-08, -3.350971e-08, -2.94404e-08, 
    1.257091e-07, -1.186311e-07, -1.058601e-08, -5.80377e-09, 2.371427e-08, 
    2.423457e-08, -7.166832e-09, -1.889276e-08, -4.807899e-09, -3.922025e-09, 
    2.326357e-08, 2.742514e-08, 3.033506e-08, -2.2905e-08, 4.965557e-09, 
    2.340985e-07, 4.407599e-08, 2.827045e-08, 2.613836e-07, 2.53611e-07, 
    1.059897e-08, -6.090792e-08, -4.376716e-09, -3.39622e-07, -2.201801e-08, 
    -1.619336e-07, -1.63413e-07, 9.164961e-08, 4.28787e-09, -1.71908e-08, 
    1.172538e-08, -2.111308e-08, 7.964474e-11, 1.985093e-09, 1.112488e-08, 
    -8.783257e-08, -5.720898e-08, 1.387036e-09, 6.97143e-08, 4.179691e-08, 
    -1.094293e-09, -1.285372e-08, -1.375821e-08, -1.957119e-10, 
    -5.152117e-09, -2.794877e-09, 6.52058e-09, -1.071104e-09, 1.156124e-10, 
    1.370807e-08,
  1.594896e-08, -1.197691e-10, -1.120213e-09, -1.514479e-09, 7.467008e-09, 
    3.963788e-08, 4.077384e-08, 7.699447e-08, 2.13177e-08, -3.256895e-08, 
    -4.614265e-09, -1.809275e-08, -6.915968e-09, -1.01465e-07, 5.974749e-08, 
    -6.709995e-08, -2.966146e-09, 8.742103e-08, 7.063164e-09, -1.848265e-07, 
    1.298514e-08, -1.554616e-08, 5.596178e-09, 1.125329e-09, -2.440487e-08, 
    -1.115927e-07, -6.053085e-09, -4.75319e-09, -6.573913e-08, -2.277483e-08, 
    -1.267414e-07, 5.895009e-08, -1.755546e-08, 1.827004e-09, 4.519489e-08, 
    -6.621912e-08, 1.624122e-08, 1.865203e-09, -1.237331e-07, 3.644902e-09, 
    8.082418e-09, 1.248719e-08, -9.605634e-08, -3.436113e-08, -3.785766e-08, 
    -2.862038e-08, -8.389549e-08, 2.722265e-08, -8.166592e-08, -1.667289e-08, 
    2.832894e-08, -6.40502e-08, -2.118518e-07, 2.207764e-09, -2.795247e-09, 
    -4.631033e-10, -1.403322e-07, -3.120603e-08, 3.642023e-08, 2.99127e-07, 
    3.470291e-10, 5.939285e-09, 5.189725e-07, -6.069899e-08, 3.47699e-08, 
    -2.209998e-08, -4.02851e-08, -6.777725e-09, -3.721669e-08, -3.52922e-08, 
    -2.055976e-07, -1.872342e-07, 1.379027e-08, -5.851405e-09, 1.193999e-08, 
    2.656208e-08, -1.73296e-08, -1.336105e-08, -4.275085e-09, -2.180553e-08, 
    2.67392e-08, 6.149453e-08, 2.866301e-08, -4.764382e-08, -2.146743e-08, 
    1.767845e-07, 8.762987e-08, 2.451367e-08, 2.651602e-07, 2.842083e-07, 
    1.659629e-08, -5.704682e-08, -5.488289e-09, -3.152766e-07, -6.086833e-08, 
    -4.864314e-07, -1.497006e-07, 2.499405e-10, 1.885934e-08, -8.644872e-09, 
    1.282393e-08, -6.020983e-09, 1.811914e-08, 9.987247e-10, 3.784777e-08, 
    -8.579372e-08, 5.998402e-09, 1.901441e-08, 6.375359e-08, 2.880762e-08, 
    -1.406022e-09, -1.482289e-08, -1.036022e-08, 5.307868e-09, -4.987612e-09, 
    -3.761454e-09, 7.725106e-09, -9.115126e-10, 8.546408e-11, 7.622134e-10,
  2.404465e-08, -4.080221e-10, -8.745928e-10, 5.142169e-09, 3.102184e-08, 
    4.166407e-08, 4.459901e-08, 6.373273e-08, 3.64995e-08, -3.282423e-08, 
    -4.171795e-08, 1.364634e-07, -9.710106e-09, -1.30845e-07, 5.602203e-08, 
    -5.249596e-08, -3.573734e-08, 2.629042e-08, -1.768387e-08, -1.195145e-07, 
    6.637606e-09, 3.812048e-07, 7.346227e-08, -7.649987e-10, -1.078649e-08, 
    -2.151512e-08, -5.848619e-09, -7.048698e-09, -7.035294e-08, 
    -1.246997e-08, -1.438497e-07, 1.303212e-07, -1.091792e-08, -3.234049e-09, 
    5.385698e-08, -6.366156e-08, 1.637407e-08, 8.242296e-11, -1.261266e-07, 
    -1.197281e-09, 2.236363e-08, 1.949104e-08, -1.995583e-07, -3.4959e-08, 
    -3.417097e-08, 7.109861e-09, -9.424002e-08, 2.323748e-08, -5.526129e-08, 
    -1.239438e-08, 2.42504e-08, -1.082764e-07, -1.994228e-07, 5.076868e-09, 
    -5.089828e-09, -2.356728e-10, -1.584509e-07, -1.320898e-08, 4.755452e-09, 
    3.922423e-07, -2.204956e-09, -8.617656e-08, 1.57048e-07, -4.480201e-08, 
    1.063716e-08, -2.339982e-08, -1.915748e-08, -3.005186e-08, -3.240677e-08, 
    -3.837579e-08, -3.020569e-07, -1.521361e-07, 1.560682e-08, 5.071684e-09, 
    -7.436256e-10, 1.3658e-08, -1.365109e-08, -7.569213e-09, -4.392035e-09, 
    -3.059688e-08, 2.678178e-08, 1.024919e-07, 2.322133e-08, -5.425966e-08, 
    -3.433786e-08, 3.422804e-08, 7.261644e-08, 4.223295e-08, 2.524232e-07, 
    2.955102e-07, 9.658493e-09, -6.696217e-08, -4.579817e-09, -2.666433e-07, 
    -6.001562e-08, -6.540454e-07, -1.460525e-07, -4.098297e-09, 3.713046e-08, 
    -6.221012e-09, 3.801449e-08, 5.594785e-09, 3.032315e-08, -1.061906e-09, 
    7.715255e-08, -5.56671e-08, 4.137121e-08, 2.244326e-08, 4.576407e-08, 
    1.14386e-08, -2.876163e-09, -5.153311e-09, 7.975245e-09, 6.003461e-09, 
    -2.492584e-09, -4.108005e-09, 8.147396e-09, -1.025462e-09, 7.506173e-11, 
    6.965968e-08,
  2.327141e-08, 1.649084e-09, 4.233129e-10, 7.267033e-09, 4.723273e-08, 
    5.235091e-08, 3.534291e-08, 5.273904e-08, 4.784164e-08, -2.726398e-08, 
    -1.605764e-08, 8.342312e-08, 9.551002e-09, -4.437726e-08, -1.52437e-09, 
    -2.03661e-08, -6.387889e-08, -1.036591e-08, 1.061602e-08, 3.506028e-08, 
    3.087604e-07, 1.081607e-07, 1.182422e-07, -2.360087e-07, -7.673009e-09, 
    -8.41402e-09, -1.723589e-08, -1.087921e-08, -8.50992e-08, -1.530844e-08, 
    -9.317392e-08, 1.489049e-07, -1.626046e-08, -1.363338e-08, 4.482757e-08, 
    -8.076182e-08, 1.509337e-08, -4.199023e-10, -1.195597e-07, -2.192736e-08, 
    3.214618e-07, 6.908351e-07, -5.903786e-08, -4.874765e-08, -2.988196e-08, 
    2.239875e-08, 1.735231e-08, 3.119652e-08, -5.146163e-08, -5.616172e-09, 
    2.030646e-08, -1.80877e-07, -1.733067e-07, 1.041966e-08, -9.740262e-09, 
    -1.129479e-10, -1.897786e-07, -3.477477e-08, -1.106845e-08, 4.175101e-07, 
    -2.367926e-09, -1.984316e-07, 7.980378e-08, -2.020716e-08, -9.418827e-09, 
    -2.470944e-08, 1.6412e-08, -4.316695e-08, -1.940413e-08, -2.595272e-08, 
    -2.59762e-07, -9.827437e-08, 2.310111e-08, -7.313304e-09, -1.757859e-08, 
    4.797073e-09, -3.873708e-09, -8.785207e-09, -5.289422e-09, 1.46543e-07, 
    2.584653e-08, 1.358219e-07, 1.373832e-08, -2.140325e-09, -3.967153e-08, 
    -6.437386e-08, 1.397452e-07, 5.529904e-08, 2.526101e-07, 2.988958e-07, 
    -1.813135e-09, -7.620248e-08, -5.66564e-09, -2.16292e-07, -2.63272e-08, 
    -6.567724e-07, -9.740162e-08, -6.404281e-08, 5.975693e-08, -1.335339e-08, 
    2.79494e-07, 1.436042e-08, 3.145792e-08, 9.713403e-10, 2.058772e-08, 
    -5.813359e-08, 6.510788e-09, 1.789948e-08, 2.204951e-08, -1.075847e-08, 
    2.526747e-09, 2.390095e-09, 1.149164e-08, -1.672862e-08, -2.072795e-09, 
    -2.955528e-09, 8.241756e-09, -1.094563e-09, 4.77911e-11, -3.645368e-10,
  1.347007e-08, 7.014705e-09, 4.339768e-09, 1.422109e-09, 1.826379e-08, 
    3.578805e-08, 2.611125e-08, 4.204969e-08, 5.555489e-08, -1.600279e-08, 
    1.232576e-07, 1.570453e-07, 4.430058e-08, -1.355068e-08, -1.435236e-07, 
    2.147853e-08, -7.447068e-08, -1.797679e-08, 1.143178e-08, 5.275467e-08, 
    1.683964e-08, -1.43387e-07, 7.830374e-08, -1.470843e-07, -3.917182e-08, 
    -6.494133e-08, -4.556375e-08, -1.711021e-08, -1.05313e-07, -1.256501e-08, 
    -7.055417e-08, 1.362831e-07, -4.795595e-08, 5.593847e-09, 4.058404e-08, 
    -1.095167e-07, 8.71363e-09, 4.15227e-10, -9.861799e-08, -6.399046e-08, 
    4.683633e-07, 8.700329e-08, 7.842877e-08, -6.351789e-08, -2.547574e-08, 
    1.080332e-08, 6.206199e-08, 3.439189e-08, -3.343546e-08, -8.240875e-11, 
    1.658731e-08, -1.397041e-07, -1.240467e-07, 1.037076e-08, -1.31144e-08, 
    -3.509513e-10, -2.056651e-07, -8.80317e-08, 2.207283e-08, 3.6724e-07, 
    -2.772367e-09, -1.267315e-07, -3.88336e-08, 2.437297e-08, -3.468163e-08, 
    -2.381773e-08, -6.284165e-08, -5.074935e-08, -8.200345e-09, 
    -8.417373e-10, -8.631605e-08, -1.082888e-07, 1.420744e-09, -4.260119e-08, 
    -8.601778e-08, -3.578862e-10, -1.33582e-12, 3.651991e-09, -4.139008e-09, 
    2.401512e-07, 2.637466e-08, 1.660536e-07, 8.784582e-10, -1.687067e-08, 
    -2.125444e-08, 5.807306e-08, 1.090694e-07, 2.596914e-08, 2.698617e-07, 
    2.915919e-07, -4.191122e-08, -8.234658e-08, -9.393631e-09, -1.108299e-07, 
    -2.520312e-08, -5.811139e-07, -9.719086e-08, -7.996982e-08, 7.693802e-08, 
    7.169568e-09, 1.780786e-07, 1.053326e-08, 2.352601e-08, 9.674018e-09, 
    -2.171987e-09, -4.31836e-08, -7.63788e-08, -7.849962e-09, -3.978698e-09, 
    -2.943011e-08, 7.890401e-08, 4.430012e-08, 6.405912e-09, -3.730304e-08, 
    -2.429488e-09, -1.662659e-09, 8.641322e-09, -1.332882e-09, -4.723049e-10, 
    -1.075231e-07,
  6.162907e-09, 2.2454e-08, 1.242796e-08, -1.074574e-08, -9.514054e-09, 
    3.480807e-09, 1.18452e-08, 2.401561e-08, 4.672751e-08, 6.235877e-08, 
    1.787961e-07, 3.783879e-08, 2.68878e-07, -1.201653e-08, -2.181792e-07, 
    4.330509e-08, -8.057985e-08, -7.601273e-09, 1.792833e-08, -7.114352e-09, 
    -1.47906e-07, -7.093269e-08, 5.527085e-08, -3.008955e-08, -1.246611e-07, 
    -1.203285e-07, -4.907048e-08, -2.047346e-08, -1.107854e-07, 
    -2.486019e-08, -7.291266e-08, 8.215756e-08, -5.300132e-08, 2.743434e-09, 
    1.395014e-07, -1.565866e-07, -9.133612e-09, 1.183196e-09, -8.71583e-08, 
    -8.61768e-08, 1.066859e-07, -2.763623e-07, 2.356614e-08, -7.262312e-08, 
    -1.674545e-08, -2.041025e-08, 4.688894e-08, -5.03826e-09, -3.056908e-08, 
    2.637364e-09, 1.279361e-08, -1.446518e-07, -7.671539e-08, 1.293955e-08, 
    -1.606007e-08, -5.840832e-09, -1.623262e-07, -1.457577e-07, 7.200759e-08, 
    2.987613e-07, -2.062848e-10, -8.41074e-08, -7.975751e-08, 7.678616e-08, 
    -4.244294e-08, -1.950372e-08, -4.258214e-08, -5.692669e-08, 
    -5.542745e-09, 1.710845e-08, 1.695156e-08, -1.200752e-07, -7.235036e-08, 
    -6.758984e-08, -2.686664e-08, -1.388173e-09, -1.194547e-08, 
    -8.045618e-09, -8.592195e-09, 5.506735e-08, 1.997734e-08, 1.908098e-07, 
    -1.599363e-08, -1.058912e-07, -4.781953e-09, -4.621654e-09, 6.186309e-08, 
    -9.495182e-09, 2.308344e-07, 2.707692e-07, 3.245731e-08, -8.427956e-08, 
    -5.858737e-09, -1.704304e-08, -4.164627e-08, -5.049026e-07, 
    -1.824482e-07, -3.521615e-08, 8.154342e-08, 9.372083e-08, -1.113761e-07, 
    2.174194e-08, 1.42345e-08, 1.871365e-08, 4.120636e-09, -3.927255e-09, 
    -9.382808e-08, -2.417602e-08, -2.74436e-08, -4.038162e-08, 4.939028e-08, 
    2.518368e-07, 6.421232e-08, 1.493788e-09, 4.34278e-09, -7.347239e-10, 
    8.734077e-09, -1.044446e-08, -9.039098e-10, -7.696968e-08,
  4.076412e-09, 5.526812e-08, 1.873622e-08, -2.043413e-08, -1.557072e-08, 
    -1.076199e-08, -9.228501e-08, -4.955194e-08, 2.964128e-08, 1.269792e-07, 
    -3.526139e-08, -1.08858e-08, 5.131325e-07, -2.060379e-07, -1.202597e-07, 
    5.600985e-08, -9.524449e-08, 2.06216e-08, 1.962078e-08, -1.194283e-07, 
    -5.74434e-08, -2.678195e-08, -5.747495e-09, 1.107622e-08, -5.953837e-09, 
    -1.557157e-07, -4.102054e-08, -1.451139e-08, -8.789465e-08, 
    -3.767747e-08, -1.20769e-08, 3.772999e-08, -5.933788e-08, -5.149843e-09, 
    3.11878e-07, -1.820335e-07, -3.652266e-08, 2.010111e-09, -7.602165e-08, 
    -8.480885e-08, -9.701513e-08, -1.181028e-07, -6.006798e-08, 
    -7.787929e-08, -1.394966e-08, -3.536087e-08, 3.559643e-08, -5.236811e-08, 
    -2.802657e-08, 4.792611e-09, 9.807835e-09, -1.841323e-07, -3.939275e-08, 
    1.778257e-08, -2.089129e-08, -3.449713e-09, -7.225259e-08, -1.951714e-07, 
    8.699099e-08, 2.09992e-07, 2.729905e-09, 4.283407e-08, -1.249122e-07, 
    1.541346e-07, -4.101861e-08, -1.294615e-08, -1.02994e-08, -5.841338e-08, 
    -9.343637e-09, 2.514543e-08, 9.23506e-08, -7.793705e-08, -1.339294e-07, 
    -5.964176e-08, 3.921414e-08, -9.923156e-10, 1.184924e-08, -2.387878e-09, 
    8.076194e-09, 1.186239e-07, 5.784102e-09, 1.974619e-07, -7.232984e-09, 
    -5.696114e-08, 2.198448e-08, -5.537282e-08, 6.896636e-08, -1.067048e-08, 
    1.861604e-07, 2.369217e-07, -3.420894e-09, -8.306461e-08, -3.230269e-09, 
    4.851034e-08, -2.535728e-09, -4.640837e-07, -2.546667e-07, 5.477688e-08, 
    7.335615e-08, 8.982906e-08, -2.08467e-08, 1.859101e-07, 5.893384e-09, 
    2.165777e-08, 1.848861e-08, 3.310248e-08, -9.691308e-08, -3.158317e-08, 
    -4.507962e-08, -4.239604e-08, 1.919062e-08, 2.49392e-08, 1.568303e-07, 
    9.673926e-08, -9.178791e-09, 2.116962e-10, 8.755705e-09, -4.724644e-09, 
    -9.054375e-10, -8.706519e-08,
  1.365123e-08, 9.148943e-08, 1.90708e-08, -1.258849e-08, 1.08102e-08, 
    -1.093178e-07, 4.666691e-08, 4.716554e-08, 1.603824e-07, -1.736834e-08, 
    -1.572878e-07, -5.634155e-08, -5.557757e-08, -1.073717e-07, 
    -4.528368e-08, 6.214188e-08, -1.284253e-07, -2.319956e-08, 1.309672e-08, 
    -1.911486e-07, -1.880318e-08, -4.946912e-09, -9.028071e-08, 5.586742e-09, 
    8.201425e-09, -2.784258e-07, -3.261181e-08, -5.462027e-09, -6.470526e-08, 
    -4.841951e-08, 1.630934e-08, 3.302165e-08, -6.542876e-08, 1.174783e-09, 
    2.075338e-07, -1.778135e-07, -6.490514e-08, 2.832735e-09, -5.883641e-08, 
    -8.411405e-08, -9.608826e-08, 6.868191e-08, -1.049392e-07, -8.329681e-08, 
    -1.285076e-08, -2.006624e-08, -2.690996e-08, -8.301063e-08, 
    -2.642124e-08, 5.387008e-09, 8.216816e-09, -8.748071e-08, -2.109708e-08, 
    2.183725e-08, -3.014716e-08, -1.55751e-10, -1.606185e-08, -1.971837e-07, 
    5.790048e-08, 1.885268e-07, 7.643706e-08, 9.509046e-08, -1.09739e-07, 
    1.752947e-07, -3.338093e-08, -5.125401e-09, 7.242591e-09, -5.631028e-08, 
    -1.093616e-08, 1.279631e-08, 7.955936e-08, -6.177623e-08, -2.01747e-07, 
    -6.621434e-08, 4.336613e-08, 8.211032e-10, 1.705018e-08, 4.066834e-09, 
    1.09664e-08, 4.099439e-08, 5.144898e-10, 1.769721e-07, -2.574455e-08, 
    2.383223e-08, 4.165287e-08, -5.536748e-08, 1.090177e-07, -4.886886e-09, 
    1.602947e-07, 1.917054e-07, -7.640409e-08, -8.757314e-08, -4.028578e-09, 
    1.026539e-07, 1.820302e-08, -4.964834e-07, -2.779437e-07, -1.386178e-08, 
    5.390035e-08, 5.75253e-08, -8.656542e-08, 2.880353e-08, -2.6156e-09, 
    2.002974e-08, 6.66883e-08, 5.67058e-08, -1.126096e-07, -3.455017e-08, 
    -5.401677e-08, -2.522478e-08, 4.881429e-09, -2.88457e-08, 2.356074e-08, 
    4.412192e-08, -3.879052e-09, 1.004185e-09, 9.046076e-09, -3.184869e-09, 
    -7.300685e-10, 2.323742e-08,
  2.859713e-08, 8.347274e-08, 2.221657e-08, 9.94828e-09, -6.490814e-08, 
    -4.551238e-07, 5.155357e-08, -4.157528e-10, -1.916158e-08, -5.37799e-08, 
    -1.226881e-07, -3.811613e-08, -1.489118e-07, -6.53331e-08, -8.309837e-08, 
    6.706467e-08, -1.509323e-07, -3.315472e-08, 1.268793e-08, -1.417748e-07, 
    -2.719651e-08, 2.203979e-08, -1.313197e-07, 8.359029e-08, -1.045884e-07, 
    -2.344992e-07, -1.87049e-08, -5.240281e-09, -5.894105e-08, -5.218772e-08, 
    -1.201784e-09, 1.720889e-08, -6.94215e-08, 5.902052e-09, 9.784844e-08, 
    -1.602964e-07, -8.548684e-08, 3.04324e-09, -3.952096e-08, -1.709526e-08, 
    -7.219833e-08, 1.071365e-07, -9.77422e-08, -8.656038e-08, -1.626984e-08, 
    2.392539e-09, -4.380257e-08, -7.353773e-08, -3.99657e-08, 3.897135e-09, 
    8.196039e-09, -9.763914e-08, -9.305233e-09, 2.289367e-08, -3.792761e-08, 
    1.399485e-10, 4.317496e-08, -1.439453e-07, -3.36403e-08, 1.537798e-07, 
    7.029348e-08, 1.150204e-08, 1.184607e-07, 1.549111e-07, 1.850348e-08, 
    -4.742674e-09, 1.19735e-09, -5.311381e-08, -1.545311e-08, 2.447678e-10, 
    4.96309e-08, -7.015512e-08, -1.912507e-07, -1.081224e-07, 3.323729e-08, 
    2.679599e-09, 2.881521e-08, -4.27471e-09, -1.929087e-08, 4.45699e-08, 
    4.634444e-09, 1.848126e-07, -5.124656e-08, 6.516541e-08, 7.974711e-08, 
    1.776834e-08, 8.819393e-08, -3.292371e-09, 1.652247e-07, 1.366881e-07, 
    1.565934e-08, -7.526978e-08, -1.308479e-09, 1.331656e-07, -9.849259e-09, 
    -5.282797e-07, -2.649893e-07, -1.111357e-08, 5.508741e-08, 1.379503e-08, 
    2.651279e-08, -1.75764e-08, 5.018713e-08, 1.49292e-08, 1.280011e-08, 
    6.128062e-08, -1.372831e-07, 9.936116e-09, -5.770323e-08, 5.929905e-10, 
    -5.820993e-09, -4.191918e-08, -2.786214e-08, -9.833911e-11, 5.551556e-09, 
    2.32169e-09, 1.15684e-08, -2.733152e-09, -5.332055e-10, 8.131894e-08,
  6.452768e-07, 6.171473e-08, 5.848079e-08, -1.384132e-08, -3.133831e-07, 
    -6.475051e-08, -3.049252e-09, -1.916607e-08, -9.129002e-08, 
    -3.908616e-08, -9.05606e-08, -5.912733e-08, -1.375499e-07, -8.905891e-08, 
    -8.717058e-08, 7.676995e-08, -1.597432e-07, 2.150301e-08, 8.164051e-09, 
    -7.519151e-08, -2.508858e-08, 5.669887e-08, -1.6702e-07, 1.901242e-09, 
    -5.322801e-08, -4.234693e-08, -2.913345e-08, -9.669634e-10, -7.65877e-08, 
    -4.686177e-08, -5.861608e-08, 7.273815e-08, -2.542919e-08, 6.069115e-09, 
    1.840567e-07, -1.625093e-07, -9.547998e-08, 2.629449e-09, -2.980806e-08, 
    1.00232e-07, -1.694849e-08, -3.113172e-08, -3.067524e-08, -8.579256e-08, 
    -1.266784e-08, 1.076859e-08, -5.842827e-08, -8.837753e-08, -1.907796e-08, 
    2.104038e-09, 7.515823e-09, -1.217983e-07, 1.52777e-08, 2.939142e-08, 
    -3.282487e-08, -4.924914e-10, 1.462837e-08, -1.187558e-07, -5.095265e-08, 
    1.215324e-07, 9.088336e-08, 3.75955e-08, -8.850208e-08, 1.451014e-07, 
    5.286083e-10, -5.791378e-09, -1.090388e-08, -4.899465e-08, -2.60041e-08, 
    -1.156951e-08, 1.815664e-08, -8.454134e-08, -9.253068e-08, -8.278204e-08, 
    9.681685e-09, 7.599397e-10, 7.947264e-09, -7.867328e-09, -1.913287e-08, 
    3.589611e-08, -8.9031e-09, 1.788192e-07, -3.619823e-08, -3.311044e-08, 
    1.491764e-07, -6.382322e-09, -5.518808e-08, 2.777938e-10, 1.721741e-07, 
    6.752208e-08, 2.234998e-08, -6.849517e-08, 5.892105e-10, 1.398787e-07, 
    -1.188738e-08, -5.307616e-07, -2.414485e-07, -2.167013e-08, 6.974011e-08, 
    -1.080167e-08, -2.117457e-08, -2.227342e-08, 1.50061e-07, 1.238692e-08, 
    -3.008893e-09, 5.709359e-08, -1.435621e-07, 1.624076e-07, 8.323872e-08, 
    2.111375e-08, -1.263078e-08, -4.737313e-08, -4.239138e-08, -5.547975e-09, 
    7.992128e-09, 3.723688e-09, 3.674117e-09, -2.723173e-09, -3.183729e-10, 
    5.038049e-08,
  9.047933e-07, 1.665115e-07, 3.701688e-07, -1.453916e-07, -1.583505e-07, 
    5.514539e-08, -1.273645e-08, -2.810771e-08, -6.406856e-08, -3.065691e-08, 
    -7.211543e-08, -5.039874e-08, -1.762903e-07, -6.836092e-08, 
    -9.632811e-08, 1.183196e-07, -1.310548e-07, 3.78098e-08, 1.449774e-08, 
    -5.7428e-08, -9.736436e-08, 7.762776e-08, -4.923629e-08, -9.897576e-10, 
    -1.998274e-09, 2.115539e-07, -3.92281e-08, -2.166871e-08, -5.682512e-08, 
    9.192263e-09, -4.499543e-08, 1.212663e-08, -5.835204e-09, 5.180482e-09, 
    1.709815e-07, -1.637412e-07, -7.934389e-08, 1.760625e-09, -2.580612e-08, 
    9.590053e-08, 4.827893e-08, 1.730391e-07, 6.105955e-08, -8.077311e-08, 
    -1.551177e-08, -3.001753e-08, -5.693511e-08, -5.838589e-08, 
    -2.024265e-08, 1.153815e-09, 7.06261e-09, -1.252565e-07, 5.721712e-08, 
    2.359643e-08, -3.027147e-08, -3.395144e-09, 4.051492e-08, -1.025056e-07, 
    -5.534876e-08, 1.083369e-07, -7.34758e-10, 3.658511e-08, -2.289324e-07, 
    1.443652e-07, 6.986348e-09, -7.229119e-09, -2.59954e-08, -4.691208e-08, 
    -4.036792e-08, -2.566458e-08, 6.52085e-09, -9.985138e-08, -1.662136e-08, 
    5.545633e-08, 7.897235e-09, -3.458467e-09, -8.370819e-09, -7.217579e-09, 
    -1.440772e-08, 6.471907e-08, -2.626763e-08, 1.563992e-07, -8.481436e-09, 
    -5.824165e-08, 9.073926e-08, 1.908472e-08, -2.395283e-07, 1.528895e-08, 
    1.177504e-07, 4.451124e-09, 1.05377e-07, -4.432388e-08, 2.698073e-10, 
    1.292287e-07, 5.072741e-08, -4.53997e-07, -2.122475e-07, -4.281594e-08, 
    6.757125e-08, -2.110266e-08, -5.447328e-08, -4.428017e-09, 4.438603e-08, 
    1.153965e-08, 4.688638e-08, 7.01632e-08, -1.019242e-07, 1.949865e-07, 
    1.757766e-07, 4.194999e-08, -2.029617e-08, -5.257425e-08, -4.778735e-08, 
    -7.29392e-09, 8.621896e-09, 4.544734e-09, 4.239737e-09, -2.457369e-09, 
    -1.934737e-10, -4.730487e-08,
  4.820333e-07, 5.422025e-07, 5.276515e-07, -4.078339e-08, 3.186813e-09, 
    6.525573e-08, -5.409794e-08, -6.07468e-08, -8.964713e-08, -3.194651e-08, 
    -4.41126e-08, -1.616155e-08, -5.382197e-07, -1.514087e-08, -7.572186e-08, 
    1.572421e-07, -1.245056e-07, 1.135396e-08, 2.379232e-08, -5.871522e-08, 
    5.559457e-09, 7.066717e-09, 1.039319e-08, -2.470244e-09, 2.171799e-08, 
    -1.682002e-08, -2.826442e-08, -2.537632e-08, -2.591997e-08, 1.912383e-09, 
    2.627661e-08, -8.30085e-08, 7.031019e-09, -3.042771e-09, -1.237964e-07, 
    -1.321169e-07, -3.438778e-08, 1.001126e-09, -2.696862e-08, 2.381518e-08, 
    7.846496e-08, -2.205581e-09, -2.183964e-08, -2.753275e-08, -3.532119e-08, 
    -5.567523e-08, -5.780993e-08, -2.733282e-08, -3.460019e-08, 2.147061e-09, 
    6.857505e-09, -3.400311e-08, 9.922707e-08, 1.817811e-08, -2.574961e-08, 
    -1.765613e-09, 3.868894e-08, -6.063725e-08, -5.711476e-08, 9.191513e-08, 
    -2.479948e-08, -2.891949e-08, -1.47426e-07, 1.334907e-07, 3.017798e-08, 
    -9.186181e-09, -3.391716e-08, -6.045804e-08, -4.484906e-08, 
    -4.503528e-08, 1.773714e-08, -9.416027e-08, -8.922308e-08, 6.590693e-08, 
    7.861956e-09, 5.828895e-09, -3.868027e-08, -4.03594e-09, -2.586481e-08, 
    9.019635e-08, -4.074064e-08, 1.468624e-07, 6.578489e-10, -5.676549e-08, 
    1.109123e-08, 8.061932e-09, -7.41673e-08, 2.614041e-08, 5.80618e-08, 
    -1.159384e-08, 4.076242e-10, -6.15195e-08, 4.199023e-10, 1.120296e-07, 
    -3.478323e-08, -2.784683e-07, -1.8704e-07, -4.41774e-08, 8.851265e-08, 
    -3.155834e-08, -2.598478e-08, 6.611174e-10, 6.801031e-08, 4.277368e-09, 
    5.711826e-08, 8.802607e-08, -8.213061e-08, 8.624755e-08, 7.467946e-08, 
    2.946894e-08, -4.827945e-08, -5.375301e-08, -4.893769e-08, -7.898109e-09, 
    1.55398e-08, 6.055291e-09, 6.617881e-09, -1.973468e-09, -4.280167e-10, 
    8.226442e-08,
  9.641496e-09, 4.301404e-08, -6.163589e-09, -1.759673e-08, 9.017964e-08, 
    3.780229e-08, -2.286221e-07, -4.748432e-08, -1.632606e-08, -1.186038e-09, 
    -3.786641e-08, 6.642955e-08, -5.979683e-08, 4.064128e-08, 1.053309e-10, 
    1.789192e-07, -1.01187e-07, -1.539479e-08, 7.380174e-08, 3.222641e-08, 
    6.448488e-09, 6.557514e-09, 4.876637e-08, -3.02299e-09, 3.097267e-08, 
    -4.012469e-08, -4.071472e-08, -1.606799e-08, -3.269946e-08, -3.01406e-08, 
    2.891358e-08, -8.39147e-08, 1.712833e-07, 1.757832e-08, -6.40909e-08, 
    -9.642855e-08, -1.237531e-08, 1.69139e-09, -5.178885e-08, -8.692075e-09, 
    5.358173e-08, -4.817451e-08, -6.807898e-08, -4.947568e-09, -2.04879e-08, 
    -7.199804e-08, -5.727361e-08, -8.599264e-08, -3.772619e-08, 3.554199e-09, 
    6.637777e-09, 1.584857e-08, 1.309779e-07, 2.368785e-08, -2.218639e-08, 
    -1.210651e-09, 2.272192e-07, -6.110157e-08, -5.804323e-08, 1.048007e-07, 
    -3.380131e-08, -4.069688e-08, -2.053895e-08, 1.141115e-07, 2.609432e-08, 
    -2.437156e-08, -3.307258e-08, -7.682257e-08, -1.903317e-08, -5.15077e-08, 
    1.851009e-08, -1.051855e-07, -1.161948e-07, -8.738709e-09, 8.306614e-09, 
    2.726779e-10, -3.913485e-08, -1.427802e-08, -2.31257e-08, -1.193126e-08, 
    -3.901238e-08, 1.299197e-07, 1.842403e-08, -1.427128e-08, 1.443135e-08, 
    1.363897e-07, -4.835221e-08, -4.089372e-09, 3.446683e-08, -2.819002e-08, 
    -3.081311e-09, -6.245047e-08, -9.506067e-09, 1.010823e-07, -6.80381e-08, 
    -1.571296e-07, -1.431699e-07, -5.457537e-10, 1.05765e-07, -3.556125e-08, 
    1.00784e-08, -3.262386e-10, -1.270207e-08, 3.982024e-09, 1.674244e-07, 
    1.187621e-07, -4.658926e-08, 1.427799e-08, -3.950839e-08, -2.541191e-08, 
    -6.558395e-08, -5.503972e-08, -5.041142e-08, -8.246786e-09, 2.410951e-08, 
    6.707341e-09, 5.016872e-09, -1.670657e-09, -6.012826e-10, -9.12911e-09,
  -2.297471e-07, -5.509969e-08, -3.596404e-08, -2.390777e-08, -1.597766e-08, 
    3.410639e-08, -1.001215e-07, -8.623033e-09, -1.525223e-09, 1.504498e-08, 
    -1.641797e-08, -1.717729e-08, 1.594424e-08, 4.582637e-08, 8.890765e-09, 
    1.939517e-07, -6.731621e-08, -2.899748e-08, 1.16465e-07, -1.940055e-08, 
    8.10212e-09, 7.368158e-09, 5.587083e-08, -3.832724e-09, 3.094647e-08, 
    -4.685535e-08, -4.430035e-09, -6.589846e-08, 6.942116e-08, -5.16211e-08, 
    5.372658e-08, -2.570749e-07, 1.764885e-07, 8.806978e-09, -4.253934e-08, 
    -5.192305e-08, -8.156245e-09, 2.797492e-09, -4.685148e-09, -2.334297e-08, 
    6.377803e-08, -6.283187e-08, -8.399047e-08, -1.97333e-08, 1.829881e-08, 
    -8.316999e-08, -5.719687e-08, -9.123883e-08, -3.486671e-08, 4.076881e-09, 
    6.482168e-09, 1.725698e-08, 1.493043e-07, 2.753791e-08, -1.97148e-08, 
    -3.546461e-10, 2.799915e-07, -9.768044e-08, -5.853381e-08, 6.515327e-08, 
    -3.855189e-08, -4.386027e-08, 6.138976e-09, 7.339381e-08, -1.691754e-08, 
    -5.792981e-08, 4.525305e-09, -7.308984e-08, 8.081884e-09, -3.360958e-08, 
    1.091166e-08, -3.593311e-08, -2.95563e-08, -4.802928e-09, 7.77834e-09, 
    -3.21379e-08, -2.87086e-08, -1.136561e-08, -1.331496e-08, -1.142314e-08, 
    -2.837555e-08, 1.2307e-07, 4.24601e-08, 2.690126e-08, 1.060812e-09, 
    9.543555e-08, -1.290044e-07, -4.457297e-08, 2.695639e-08, -3.986969e-08, 
    -4.59147e-09, -5.316287e-08, -1.010349e-08, 8.845706e-08, 1.125833e-07, 
    -2.520411e-07, -1.041518e-07, 9.734356e-08, 1.055004e-07, -4.359515e-08, 
    1.14843e-07, -8.894929e-10, -3.514376e-08, 3.064329e-09, 1.340708e-07, 
    7.69802e-08, 5.212996e-08, -1.537296e-08, -6.348785e-08, -5.138577e-08, 
    -8.405823e-08, -5.703487e-08, -5.094091e-08, -8.443862e-09, 2.374679e-08, 
    9.434848e-09, 1.266386e-09, -3.318323e-09, -6.158842e-10, 1.118678e-09,
  -2.582457e-07, -5.881537e-08, -4.225916e-08, -2.404335e-08, -3.399276e-08, 
    -2.976134e-08, -3.074905e-08, -9.863868e-09, 4.400192e-09, 1.009317e-08, 
    -7.321148e-09, -1.925531e-08, 1.358927e-08, 3.991823e-08, 1.126506e-08, 
    2.121442e-07, -4.482346e-08, 3.122005e-08, 1.018677e-07, -1.839425e-08, 
    8.011568e-09, 4.274909e-09, 5.868748e-08, -4.979199e-09, 3.443535e-08, 
    -4.887914e-08, -6.305243e-09, -1.568441e-08, 1.967274e-07, -2.361621e-07, 
    -1.170832e-08, 1.607606e-08, 3.818997e-08, -1.655451e-09, -1.116695e-08, 
    7.332631e-09, -4.964829e-09, 3.395456e-09, 3.134035e-07, -3.050224e-08, 
    7.141985e-08, -6.563226e-08, -8.892948e-08, -1.11641e-08, -6.164959e-08, 
    -6.743988e-08, -5.749058e-08, -9.972172e-08, -3.314329e-08, 3.774716e-09, 
    6.312433e-09, 1.628069e-08, 1.558912e-07, 2.81707e-08, -1.815673e-08, 
    -1.448939e-10, 8.688045e-08, -1.172494e-07, -5.887681e-08, 6.416136e-08, 
    -3.882968e-08, -4.352472e-08, 7.915446e-10, 7.491737e-08, -2.135529e-08, 
    -4.453585e-08, -1.402458e-08, -3.737966e-09, -4.421207e-08, 
    -1.583447e-08, 1.570982e-09, 3.394887e-07, -1.151619e-08, -4.491028e-09, 
    7.36712e-09, -2.006499e-08, -1.763124e-08, -9.521614e-09, -9.784941e-09, 
    -1.071265e-08, 1.735827e-09, 1.197105e-07, 3.992051e-08, 2.35662e-08, 
    -2.034483e-09, 6.834836e-08, -1.719238e-07, -3.950021e-08, 1.68287e-08, 
    -3.829388e-08, -5.250683e-09, -5.055316e-08, -9.490179e-09, 8.708604e-08, 
    1.055838e-07, -3.272328e-07, -1.017089e-07, 8.653643e-08, 1.040551e-07, 
    -2.043602e-08, 6.374427e-08, -5.820482e-10, -5.190256e-08, 2.357439e-09, 
    4.923874e-08, 1.17596e-08, 1.602314e-07, -2.330029e-08, -7.070906e-08, 
    -6.42562e-08, -9.977583e-08, -5.853934e-08, -5.124338e-08, -8.585346e-09, 
    1.278573e-08, 3.924981e-09, 6.755982e-09, -1.897448e-09, -8.982681e-11, 
    -5.429115e-10,
  -3.035052e-07, -5.994912e-08, -4.397145e-08, -2.402169e-08, -3.831872e-08, 
    -4.242781e-08, -1.80122e-08, -1.176841e-08, 6.69354e-09, 1.291744e-08, 
    -1.322064e-09, -1.026353e-08, 1.045964e-08, 3.7105e-08, 1.294507e-08, 
    2.367775e-07, -2.509316e-08, 2.800186e-08, 9.072008e-08, -1.78693e-08, 
    7.676022e-09, -9.686119e-10, 5.971469e-08, -5.400693e-09, 3.688285e-08, 
    -4.930371e-08, 4.02008e-09, -2.529998e-08, 8.974325e-09, -7.041842e-08, 
    -2.302079e-08, -3.038679e-08, 3.772425e-08, 1.306432e-08, -9.407586e-09, 
    3.825835e-08, 2.883428e-09, 3.736616e-09, 2.281843e-07, -3.108451e-08, 
    4.746974e-08, -6.852918e-08, -9.044805e-08, -1.130003e-08, -7.196149e-09, 
    -9.964037e-08, -5.7715e-08, -9.380847e-08, -3.064065e-08, 3.569326e-09, 
    6.151367e-09, 1.588262e-08, 1.575007e-07, 2.942415e-08, -1.731856e-08, 
    3.015714e-09, 4.669721e-08, -1.317035e-07, -5.907498e-08, 7.61634e-08, 
    -3.85262e-08, -4.208698e-08, 1.758849e-09, 7.731619e-08, -1.356639e-08, 
    5.052857e-08, 6.328185e-08, 3.868763e-09, 2.067509e-09, -3.863545e-08, 
    -8.084839e-09, 4.751709e-07, 7.085873e-09, -4.536673e-09, 6.486658e-09, 
    6.943196e-09, -2.242193e-08, -8.241585e-09, -4.151985e-10, -9.682594e-09, 
    -1.167763e-08, 1.171105e-07, 3.695897e-08, 2.257207e-08, -1.245439e-09, 
    7.219978e-08, -1.730773e-07, -3.729508e-08, 1.373353e-08, -3.185232e-08, 
    -5.937181e-09, -3.574003e-08, -8.77975e-09, 8.527685e-08, 1.346734e-08, 
    -3.598729e-07, -1.038606e-07, 5.157472e-08, 9.825055e-08, -1.194971e-08, 
    -1.585863e-08, -9.512888e-10, -5.396046e-08, 1.082228e-09, 4.66755e-08, 
    1.64215e-08, -1.356074e-07, -2.76093e-08, -7.438166e-08, -6.790015e-08, 
    -1.036909e-07, -5.934805e-08, -5.132677e-08, -8.718189e-09, 6.217419e-09, 
    4.258482e-09, 5.490605e-09, -1.4813e-09, 6.102141e-11, -2.215074e-09,
  -3.382739e-07, -5.974033e-08, -4.222619e-08, -2.421967e-08, -4.002203e-08, 
    -4.743919e-08, 7.472238e-09, -1.447489e-08, 7.925735e-09, 1.439474e-08, 
    5.251763e-10, -1.018674e-08, 7.605479e-09, 4.08873e-08, 1.412656e-08, 
    2.700999e-07, -1.876012e-08, 3.010183e-08, 8.50947e-08, -1.869404e-08, 
    7.311939e-09, -5.143249e-09, 5.992712e-08, -5.69986e-09, 3.763915e-08, 
    -4.956536e-08, 4.339995e-10, -4.608461e-08, -6.407788e-09, -5.419162e-08, 
    -2.085011e-08, -2.804228e-08, 3.780741e-08, 5.165305e-09, -5.156664e-09, 
    4.175791e-08, 9.899816e-09, 3.094286e-09, 1.600661e-07, -3.398944e-08, 
    4.110464e-08, -7.097952e-08, -9.163986e-08, -1.776746e-08, 1.834604e-08, 
    -1.119293e-07, -5.788917e-08, -8.953714e-08, -2.747412e-08, 5.887017e-09, 
    5.981676e-09, 1.560812e-08, 1.568053e-07, 3.086135e-08, -1.692714e-08, 
    6.249707e-09, 7.933983e-08, -1.404819e-07, -5.931185e-08, 8.143195e-08, 
    -3.763608e-08, -3.992312e-08, 2.483546e-09, 4.252755e-08, -1.111506e-08, 
    1.522511e-08, 6.1869e-08, -1.567929e-08, 1.582924e-08, -1.853499e-08, 
    -6.068547e-09, 4.915045e-07, -2.753399e-08, -4.55492e-09, 5.553453e-09, 
    -1.998734e-08, -2.527945e-08, -6.527671e-09, -1.023842e-09, 
    -8.600352e-09, -1.286276e-08, 1.142818e-07, 3.27525e-08, 2.097141e-08, 
    -1.218325e-09, 7.286252e-08, -1.613617e-07, -3.579277e-08, 1.636672e-08, 
    -2.708316e-08, -5.315371e-09, -2.46968e-08, -8.721941e-09, 8.313384e-08, 
    -2.053753e-10, -4.16273e-07, -1.11991e-07, 4.275131e-08, 9.145975e-08, 
    -1.178154e-08, -1.728273e-08, -1.918359e-09, -5.667984e-08, 
    -1.947718e-09, 4.515056e-08, 1.657378e-08, -8.723958e-08, -3.038514e-08, 
    -7.666398e-08, -6.975614e-08, -1.055396e-07, -5.974522e-08, 
    -5.138867e-08, -8.829318e-09, 4.839137e-09, -2.089871e-09, -1.07903e-09, 
    -1.048281e-09, -3.096972e-10, -3.604839e-09,
  -3.385018e-07, -6.087691e-08, -4.166145e-08, -2.398281e-08, -4.114167e-08, 
    -5.019649e-08, 7.29824e-09, -1.562705e-08, 8.841198e-09, 1.562694e-08, 
    1.501462e-09, -1.110379e-08, 4.845106e-09, 4.580124e-08, 1.647413e-08, 
    2.877614e-07, -1.63612e-08, 2.979937e-08, 8.561703e-08, -1.971455e-08, 
    4.920821e-09, -6.219238e-09, 5.973743e-08, -6.225036e-09, 3.756838e-08, 
    -5.223717e-08, -2.043294e-09, -4.489743e-08, -1.179524e-08, 
    -5.718653e-08, -1.836952e-08, -4.516028e-08, 3.668424e-08, 7.029371e-09, 
    -2.901288e-09, 4.149786e-08, 1.490537e-08, 1.239371e-09, 1.876324e-07, 
    -3.377836e-08, 2.591995e-08, -7.319977e-08, -9.302363e-08, -1.494059e-08, 
    4.620642e-08, -1.186721e-07, -5.831669e-08, -8.781959e-08, -2.382851e-08, 
    1.686665e-09, 5.786958e-09, 1.554838e-08, 1.549908e-07, 3.266982e-08, 
    -1.683429e-08, -3.444711e-10, 1.103343e-07, -1.454492e-07, -5.977719e-08, 
    8.203504e-08, -3.647881e-08, -3.927994e-08, 3.148898e-09, 2.945897e-08, 
    -1.320661e-08, -3.390539e-08, 6.890673e-08, -1.802562e-08, 2.527895e-08, 
    -1.626995e-08, -1.816261e-09, 2.817093e-07, -2.946274e-08, -4.597155e-09, 
    4.580279e-09, -2.633658e-08, -2.742179e-08, -4.913602e-09, -3.771277e-10, 
    -7.276753e-09, -9.482221e-09, 1.111003e-07, 2.972638e-08, 1.933017e-08, 
    -2.428806e-09, 7.321671e-08, -1.558996e-07, -3.497223e-08, 1.770348e-08, 
    -2.028492e-08, -4.751541e-09, -1.876676e-08, -1.055344e-08, 8.055154e-08, 
    -6.618052e-09, -4.453761e-07, -1.11621e-07, 4.30199e-08, 8.572704e-08, 
    -9.631686e-09, -1.929163e-08, -3.62963e-09, -6.033009e-08, -1.737007e-09, 
    4.401841e-08, 1.590308e-08, -7.721485e-08, -3.240712e-08, -7.83549e-08, 
    -7.095105e-08, -1.065863e-07, -5.995048e-08, -5.145637e-08, 
    -8.931238e-09, 4.39718e-09, -1.121498e-09, 2.218385e-09, 3.363922e-10, 
    -7.55648e-10, -4.225626e-09,
  -3.334942e-07, -6.025653e-08, -4.368326e-08, -2.130457e-08, -4.246738e-08, 
    -5.250251e-08, 1.050819e-08, -1.786532e-08, 9.748192e-09, 1.67239e-08, 
    2.030106e-09, -1.139517e-08, 2.711431e-09, 4.98261e-08, 1.531578e-08, 
    2.333841e-07, -1.380115e-08, 2.905432e-08, 8.529321e-08, -2.033414e-08, 
    1.605144e-09, -7.355652e-09, 5.891889e-08, -6.864866e-09, 3.692173e-08, 
    -5.412278e-08, 7.083827e-10, -4.364733e-08, -1.506805e-08, -5.176207e-08, 
    -1.611272e-08, -3.783748e-08, 3.210755e-08, 3.724949e-09, -8.75275e-10, 
    4.292747e-08, 1.845555e-08, -7.712089e-10, 1.635786e-07, -3.487747e-08, 
    5.043262e-09, -7.542462e-08, -9.376453e-08, -1.033174e-08, 5.104278e-08, 
    -1.260387e-07, -5.890308e-08, -8.604948e-08, -2.112749e-08, 2.747043e-09, 
    5.522281e-09, 1.598312e-08, 1.524984e-07, 3.107973e-08, -1.690601e-08, 
    -6.657842e-09, 1.514021e-07, -1.479086e-07, -6.05037e-08, 7.590906e-08, 
    -3.485184e-08, -3.8336e-08, 3.708124e-09, 2.164397e-08, -8.71637e-09, 
    -3.580942e-08, 6.462471e-08, -2.347133e-08, 3.205048e-08, -1.562125e-08, 
    3.309879e-09, 6.744676e-08, -3.221055e-08, -3.98245e-09, 3.456009e-09, 
    5.780976e-09, -2.828791e-08, -4.372566e-09, 9.418271e-10, -5.68366e-09, 
    -9.68646e-09, 1.071465e-07, 2.821798e-08, 1.764283e-08, -7.047674e-09, 
    7.309325e-08, -1.498209e-07, -3.340335e-08, 1.673196e-08, -1.297542e-08, 
    -5.572133e-09, -1.620156e-08, -1.165844e-08, 7.626047e-08, -9.61461e-09, 
    -4.569368e-07, -1.10949e-07, 4.057995e-08, 8.132497e-08, -8.320012e-09, 
    -1.921092e-08, -6.272465e-09, -6.199306e-08, -1.610793e-09, 4.32334e-08, 
    1.442265e-08, -6.889127e-08, -3.39503e-08, -7.969015e-08, -7.187032e-08, 
    -1.073228e-07, -6.009623e-08, -5.150628e-08, -9.040605e-09, 4.235176e-09, 
    3.801767e-09, 2.723766e-09, -1.703974e-09, -9.233716e-10, -4.165599e-09,
  -3.293956e-07, -5.615289e-08, -4.28721e-08, -1.979049e-08, -4.376113e-08, 
    -5.370941e-08, 9.71022e-09, -1.934745e-08, 1.138096e-08, 1.785554e-08, 
    2.16221e-09, -1.130365e-08, -1.635954e-10, 5.081461e-08, 1.433659e-08, 
    1.167905e-07, -1.420258e-08, 2.807576e-08, 8.364809e-08, -2.125284e-08, 
    4.234835e-10, -9.460791e-09, 5.670438e-08, -8.230586e-09, 3.544187e-08, 
    -5.354934e-08, 2.857064e-09, -3.519767e-08, -1.735191e-08, -6.508071e-08, 
    -1.319961e-08, -2.815159e-08, 2.919796e-08, -4.510866e-09, -8.599272e-10, 
    4.324261e-08, 2.143672e-08, -2.712284e-10, -1.716694e-07, -3.760591e-08, 
    -2.201574e-08, -7.68855e-08, -9.295755e-08, -7.444598e-09, 5.272648e-08, 
    -1.323165e-07, -5.942775e-08, -8.697327e-08, -1.988149e-08, 2.907029e-09, 
    5.14234e-09, 1.68551e-08, 1.490756e-07, 3.263006e-08, -1.721835e-08, 
    -6.005848e-09, 1.968069e-07, -1.498205e-07, -6.157258e-08, 7.033124e-08, 
    -3.223658e-08, -3.594084e-08, 3.138211e-09, 1.930668e-08, 3.703732e-09, 
    -3.508262e-08, 6.396056e-08, -2.750926e-08, 2.542151e-08, -1.419028e-08, 
    6.583377e-09, 1.099429e-07, -3.326102e-08, -4.242224e-09, 1.96605e-09, 
    5.702873e-09, -2.926224e-08, -3.537536e-09, 8.452584e-09, -4.606591e-09, 
    -1.052024e-08, 1.020624e-07, 3.285732e-08, 1.560363e-08, -1.111675e-08, 
    7.34351e-08, -1.45849e-07, -3.074206e-08, 1.364783e-08, -2.252307e-09, 
    -7.143399e-09, -1.625513e-08, -1.184432e-08, 7.261666e-08, -1.188687e-08, 
    -4.566917e-07, -1.079377e-07, 4.013498e-08, 7.608389e-08, -6.464825e-09, 
    -1.845569e-08, -8.993958e-09, -6.257661e-08, -1.347246e-09, 4.258084e-08, 
    1.24021e-08, -5.867548e-08, -3.518289e-08, -8.083896e-08, -7.267386e-08, 
    -1.079659e-07, -6.025607e-08, -5.153913e-08, -9.173277e-09, 4.1872e-09, 
    3.625098e-09, 6.885116e-09, -4.774385e-09, -3.022869e-09, -5.772904e-09,
  -3.255855e-07, -4.940938e-08, -3.945564e-08, -1.681502e-08, -4.587088e-08, 
    -5.788837e-08, 7.62742e-09, -1.913151e-08, 1.375139e-08, 1.972836e-08, 
    2.169315e-09, -1.056543e-08, -3.62769e-09, 4.735153e-08, 1.324059e-08, 
    3.036368e-08, -8.622919e-09, 2.780683e-08, 8.00907e-08, -2.280643e-08, 
    -3.802313e-09, -1.43479e-08, 5.005205e-08, -1.110999e-08, 3.18941e-08, 
    -5.149167e-08, 3.727621e-09, -3.211761e-08, -1.905852e-08, -7.583861e-08, 
    -7.288065e-09, -2.074665e-08, 2.219082e-08, -3.316387e-08, -3.164416e-09, 
    4.265331e-08, 2.461378e-08, -1.03681e-09, -2.971109e-07, -4.305293e-08, 
    -6.181193e-08, -7.685122e-08, -9.158927e-08, -6.635688e-09, 5.130056e-08, 
    -1.398199e-07, -5.930036e-08, -9.084496e-08, -1.990869e-08, 2.765127e-09, 
    4.483326e-09, 1.895063e-08, 1.442299e-07, 3.709741e-08, -1.776675e-08, 
    -5.896993e-09, 2.342072e-07, -1.429857e-07, -6.280645e-08, 6.823679e-08, 
    -2.696135e-08, -2.991311e-08, -3.369109e-10, 1.387001e-08, 5.804305e-08, 
    -3.376857e-08, 5.957219e-08, -2.785231e-08, 2.700148e-08, -1.222014e-08, 
    9.491202e-09, -7.591638e-08, -3.016243e-08, -3.333469e-09, -7.9757e-10, 
    -1.213886e-08, -2.768186e-08, -2.964356e-09, 7.27716e-09, -4.49387e-09, 
    -1.197566e-08, 9.369174e-08, 3.653338e-08, 1.220786e-08, -1.370819e-08, 
    7.015916e-08, -1.252811e-07, -2.494875e-08, 1.194121e-08, -2.76907e-09, 
    -1.02296e-08, -1.510524e-08, -1.101947e-08, 6.678115e-08, -1.102757e-08, 
    -4.410814e-07, -1.006045e-07, 3.414306e-08, 6.87948e-08, -4.540527e-09, 
    -1.708776e-08, -1.365016e-08, -5.922176e-08, -1.087038e-09, 4.179793e-08, 
    8.237919e-09, -3.63969e-08, -3.633903e-08, -8.218461e-08, -7.364184e-08, 
    -1.087605e-07, -6.056194e-08, -5.156556e-08, -9.414237e-09, 4.071296e-09, 
    2.574325e-10, -4.263256e-14, 2.310134e-09, -9.35276e-09, -1.454225e-09,
  -2.464214e-13, -4.958769e-13, -4.542975e-13, -2.4986e-13, 4.895363e-14, 
    1.456307e-13, -2.352739e-14, 9.143466e-14, 3.490215e-13, -2.39981e-13, 
    -5.096608e-13, 2.747745e-14, 3.391868e-13, -6.732532e-14, 7.998363e-14, 
    1.347849e-14, -3.33148e-13, 6.022345e-13, -7.817667e-14, 1.441265e-14, 
    -1.139078e-12, -1.839239e-12, -3.403585e-13, 4.282571e-13, -5.972708e-13, 
    1.946253e-14, 6.206366e-14, 3.319811e-14, 2.705117e-14, 3.695416e-14, 
    1.337228e-14, 9.10757e-14, -5.451802e-15, 1.121644e-13, 2.050182e-14, 
    -1.383342e-14, 4.620882e-13, -5.598351e-12, -4.401517e-13, 1.976138e-13, 
    2.256211e-13, -1.068791e-12, -1.397932e-13, 2.40414e-13, 1.535259e-13, 
    2.02624e-13, 8.611466e-14, 8.267809e-13, 2.838863e-12, 1.193058e-12, 
    -2.580826e-12, 1.962989e-14, 3.408214e-13, -4.194262e-13, 3.21963e-13, 
    -7.117361e-13, 3.083766e-13, -2.107382e-13, 1.497642e-13, -6.994812e-13, 
    9.772362e-13, -7.929094e-13, 1.03493e-12, -6.31642e-13, 1.547424e-13, 
    5.5754e-13, -1.078241e-13, -1.399172e-13, 2.926162e-13, 1.249223e-13, 
    -2.731107e-13, -1.674656e-13, 7.781766e-14, 2.475111e-13, -6.548424e-14, 
    1.405096e-13, -1.973944e-13, -1.856023e-12, -1.273902e-12, -3.340637e-13, 
    -7.254759e-14, 4.840393e-13, -2.485863e-14, -1.701701e-13, 4.029749e-15, 
    4.167672e-14, -4.121198e-13, 7.786137e-13, 7.221139e-13, 2.366483e-14, 
    1.470491e-13, 2.894652e-12, -1.945564e-13, 2.096338e-13, -9.574096e-14, 
    -2.428854e-13, 1.132324e-13, 3.258955e-13, 1.238385e-13, 4.714579e-13, 
    -6.97137e-13, 1.008701e-13, 8.265784e-13, 2.495295e-12, 9.943909e-14, 
    6.113679e-13, 4.895718e-13, 5.931793e-13, 8.078414e-13, 5.15059e-13, 
    3.888437e-13, -5.210287e-14, -1.694452e-15, -7.802643e-14, 4.52405e-13, 
    -1.824787e-12, 3.568946e-13, -4.83764e-13, 1.654774e-12, -1.284458e-12,
  -2.275778e-13, -2.200619e-13, -2.875999e-13, -3.648594e-13, -4.016831e-13, 
    -3.816628e-13, -4.432385e-13, -2.59845e-13, -1.512088e-13, -6.990064e-14, 
    -5.589047e-14, -1.71986e-13, 5.75876e-14, -3.018193e-13, -2.006135e-13, 
    2.895111e-13, 1.035573e-13, -2.49678e-13, -7.482758e-14, 3.048474e-13, 
    4.698469e-13, 3.887396e-13, 1.09633e-12, -6.310719e-14, 8.340645e-15, 
    -1.653486e-13, -7.472982e-13, -1.206549e-13, -3.135357e-14, 4.16024e-14, 
    2.060194e-14, 1.462696e-13, -1.360172e-13, -1.571469e-13, 7.826144e-14, 
    -1.132395e-13, 3.821679e-13, -1.362033e-13, -1.93358e-13, -4.935913e-13, 
    -1.121579e-12, 2.430211e-14, -1.055788e-13, -5.949429e-14, -1.208836e-12, 
    -1.884078e-12, -9.583918e-13, 1.748276e-13, 1.727178e-13, 8.656381e-13, 
    -7.122239e-15, -4.881959e-15, 6.558611e-13, -2.069625e-12, 2.803084e-13, 
    -5.564226e-13, -3.046627e-13, -1.135097e-12, -2.810991e-13, 
    -2.887232e-12, -3.195157e-13, -1.226526e-13, -8.657882e-14, 
    -1.956647e-14, -4.201025e-13, 1.166304e-13, 1.806164e-13, 4.065491e-14, 
    -1.730318e-13, 7.65433e-14, 8.026129e-13, 1.633726e-13, -4.001337e-13, 
    8.332212e-14, -4.303314e-15, -9.117575e-13, 5.912041e-13, 6.894532e-13, 
    -4.344935e-12, -7.286929e-13, -1.087017e-13, -9.432352e-14, -1.35224e-12, 
    8.477851e-15, -1.870337e-12, -1.209416e-12, -6.603731e-13, 3.475407e-13, 
    -1.666432e-12, -3.694674e-13, 4.814339e-14, 2.208024e-13, 1.000661e-12, 
    -1.111069e-12, -8.84437e-14, 8.206601e-13, -3.236547e-13, -6.135751e-14, 
    3.7535e-13, 4.328314e-13, -8.736757e-14, -4.876714e-15, 2.042509e-13, 
    -6.469813e-12, 7.88359e-13, 6.156871e-13, 7.737337e-13, 2.195589e-12, 
    1.413168e-12, 5.555364e-13, 3.444904e-13, -7.587531e-15, -1.651153e-13, 
    -2.615053e-13, 1.032135e-13, -4.812541e-14, -9.297591e-13, 7.270158e-12, 
    9.80103e-14, 2.742476e-15,
  6.786238e-15, -3.849698e-14, -1.245531e-13, -2.03601e-13, -1.815076e-13, 
    -4.100886e-14, 1.509765e-13, 3.835265e-13, 2.807615e-13, 1.748601e-13, 
    -9.714451e-15, -1.781214e-13, -5.320744e-14, 1.530442e-13, 4.982958e-13, 
    4.275386e-13, 9.953288e-14, 1.961695e-13, -2.171839e-13, -4.402867e-13, 
    4.345968e-13, 4.609924e-13, 3.03535e-13, -1.482564e-13, 1.054296e-13, 
    6.97456e-13, 3.418377e-13, 4.601874e-14, 4.95437e-14, 1.740275e-13, 
    -8.926193e-14, 4.997391e-14, -1.01863e-13, -7.99083e-14, 5.381806e-14, 
    1.726536e-13, -1.944743e-12, -3.823625e-13, -2.960132e-14, -1.018173e-12, 
    2.887135e-13, -1.709605e-13, -3.584251e-13, 1.140995e-13, -8.332224e-14, 
    6.824263e-13, -8.08513e-13, -6.723788e-14, -5.150963e-13, -2.261646e-14, 
    -1.502826e-13, 9.939272e-14, -5.633133e-14, -1.871792e-11, 2.761343e-13, 
    1.500446e-12, 1.564027e-13, -1.476561e-12, 1.557948e-13, 1.035307e-12, 
    8.987255e-13, -6.888379e-13, 4.496958e-13, 1.656342e-13, 4.703515e-13, 
    -4.44228e-14, 1.386391e-13, -1.207368e-15, -3.920475e-14, -3.455569e-14, 
    -1.220954e-12, 1.006278e-13, 1.12281e-12, 5.037637e-14, -5.366999e-13, 
    8.493622e-13, -5.175461e-13, 4.034932e-13, -5.484397e-12, -9.002382e-13, 
    2.793946e-13, 1.638308e-13, 6.993503e-13, 8.432144e-14, -3.979317e-13, 
    6.977752e-13, -1.72036e-12, -1.870448e-13, -2.001725e-12, -1.078047e-12, 
    -1.827566e-13, -1.085992e-13, 3.080036e-13, -1.583329e-12, 1.378758e-13, 
    2.124467e-13, -7.746609e-13, -1.31839e-13, 7.46847e-13, 1.116413e-12, 
    -2.984279e-13, -9.953757e-14, 3.917665e-13, -1.101951e-12, -1.253581e-13, 
    -1.113415e-13, -7.076284e-14, -4.710121e-13, -7.490397e-13, 
    -1.314573e-12, -1.491376e-12, -5.144773e-13, -5.868639e-13, 
    -5.919709e-13, -5.8821e-13, 1.208349e-12, 2.114735e-12, 1.869708e-11, 
    -1.044377e-12, -7.155387e-14,
  2.674666e-13, 2.889911e-13, 2.45276e-13, 1.935396e-13, 1.831313e-13, 
    2.539219e-13, 3.173573e-13, 3.946565e-13, 1.963013e-13, 3.372302e-14, 
    -7.185919e-14, -3.985146e-13, -2.977341e-13, -7.711748e-13, 
    -6.806916e-13, 2.462613e-13, 1.993725e-13, 1.963221e-13, 3.525982e-13, 
    8.151813e-14, -9.944823e-14, 1.02654e-13, 4.048845e-13, 3.636119e-13, 
    6.390583e-13, -1.002115e-13, -3.565204e-14, 9.588164e-14, 3.413242e-13, 
    5.308254e-14, -1.187522e-13, -3.358425e-14, -5.691142e-13, -5.422052e-14, 
    -3.097522e-13, -3.337053e-13, -3.023158e-12, 1.989176e-12, -1.890293e-13, 
    -5.757423e-13, 2.467859e-13, 1.571604e-12, -2.283868e-13, 7.280244e-14, 
    1.767197e-13, 6.194212e-13, -1.746152e-12, -6.889975e-13, 2.81497e-13, 
    -1.298935e-13, -9.30242e-13, 2.515765e-12, -5.408729e-13, 3.131434e-12, 
    8.995339e-14, 2.661191e-12, -3.1051e-12, -6.182193e-13, 2.264536e-13, 
    1.255166e-12, 1.918604e-13, -4.882622e-13, 9.876405e-13, 1.895872e-13, 
    6.389888e-14, 1.110737e-12, 2.176037e-14, 8.493206e-14, 1.004891e-13, 
    -3.998191e-13, -1.947054e-14, 1.039419e-12, 7.632783e-13, -4.826695e-14, 
    -8.835474e-13, 6.138146e-14, 1.102675e-12, 3.175533e-12, -1.277558e-11, 
    -1.94289e-15, 9.900344e-13, -9.62705e-13, 1.854281e-13, -8.732737e-13, 
    -1.723621e-14, -4.124617e-13, -9.172385e-13, 3.082951e-13, -1.136086e-12, 
    -8.640796e-13, -2.935291e-13, -1.400802e-12, 4.737669e-13, 7.302811e-13, 
    4.108242e-13, -1.770134e-11, -4.740152e-13, 2.957495e-13, -5.724934e-12, 
    -1.613293e-13, -1.082676e-12, -8.423028e-13, 4.00755e-13, -4.851406e-13, 
    -2.745304e-13, -7.781276e-14, 2.085832e-14, -5.765249e-13, -3.562844e-13, 
    -2.968042e-13, -9.012791e-13, -5.582618e-13, -3.342326e-13, 3.774758e-15, 
    -5.651035e-14, 1.101856e-12, -1.636923e-12, -1.374299e-12, -1.185094e-13, 
    -6.192824e-13,
  5.754147e-13, 7.665951e-13, 7.012585e-13, 6.711159e-13, 5.020012e-13, 
    1.905004e-13, 1.397632e-13, 7.518569e-13, 5.987016e-13, -4.418826e-13, 
    -4.469897e-13, -7.090023e-13, -5.592887e-13, -7.738393e-13, 4.4513e-13, 
    2.182421e-13, 1.573464e-13, 1.739719e-13, 3.786971e-13, 1.643824e-13, 
    -3.701345e-13, -6.350059e-13, -2.337158e-13, 3.754913e-13, -3.621409e-13, 
    -4.460737e-13, 5.626194e-13, 4.155704e-13, 3.040623e-14, 4.877626e-13, 
    5.494355e-13, -5.565687e-13, -3.182871e-13, -4.36734e-14, -2.904621e-14, 
    -3.869544e-13, -1.200043e-12, 7.228246e-13, 6.806361e-13, -1.169845e-12, 
    -1.026818e-13, -9.909157e-13, 1.202649e-13, -4.27075e-13, 1.250958e-12, 
    1.460568e-12, -3.778922e-14, -9.443141e-14, -6.326328e-14, 1.400289e-11, 
    7.464307e-13, 2.361569e-12, 4.918898e-13, -2.033204e-12, 4.543657e-14, 
    1.343897e-12, -9.763995e-13, -2.313113e-12, -1.65537e-13, 6.952772e-13, 
    -4.251183e-13, -8.383155e-13, -5.62092e-13, 5.959399e-14, -2.659622e-13, 
    2.786521e-13, 1.848383e-13, 3.939904e-14, 3.397976e-13, 2.212022e-12, 
    9.400397e-13, -1.185024e-13, 1.919437e-13, -4.678896e-13, -8.017948e-13, 
    5.48589e-14, -4.810492e-13, -6.728229e-13, -4.567439e-12, -4.048151e-14, 
    3.589073e-13, 1.086168e-12, 3.889528e-13, 3.110984e-13, 5.637851e-13, 
    -1.020364e-12, 1.462858e-13, 5.694195e-13, -1.221866e-12, -5.482836e-13, 
    -1.517536e-13, 8.845341e-13, 3.613845e-13, 9.991369e-13, -2.656347e-13, 
    1.051412e-11, 1.911721e-13, -2.974981e-13, -8.266998e-14, 9.395124e-13, 
    5.724449e-13, 4.760775e-13, 1.134544e-12, 8.84709e-15, -1.813688e-13, 
    -3.912565e-13, -8.330836e-14, 2.116224e-13, -7.277928e-13, -3.639172e-13, 
    -7.488871e-13, -5.982853e-13, -1.876138e-13, 2.573081e-13, 1.288553e-13, 
    1.98378e-12, 1.433311e-11, -5.831224e-12, -1.261434e-12, -7.476103e-13,
  3.63265e-13, 6.225576e-13, 9.332535e-13, 7.66387e-13, 3.472778e-13, 
    4.15723e-13, -4.710121e-13, -2.399192e-13, -4.224954e-13, -9.158785e-13, 
    7.549517e-15, 3.578249e-13, -1.253997e-13, 9.825474e-15, -7.520651e-13, 
    3.411937e-13, -4.772127e-13, -1.949274e-13, -1.416575e-13, 2.670086e-14, 
    -1.56658e-12, -2.437606e-12, -2.817468e-12, -1.827649e-12, -1.317224e-12, 
    -1.802059e-12, -9.914292e-14, 7.898682e-13, -1.389167e-12, -1.120048e-12, 
    -3.532397e-12, -4.799994e-12, -6.242784e-13, -9.237056e-14, 
    -2.067069e-12, 5.530021e-13, -7.108592e-13, -5.964257e-13, 1.933897e-12, 
    -3.921141e-13, 6.559086e-13, -2.93382e-12, 1.781492e-13, -4.56666e-13, 
    4.513112e-12, 8.030798e-13, -4.640455e-13, -2.049902e-12, -2.317857e-12, 
    1.00057e-11, 4.537551e-13, -6.439294e-15, -2.115047e-12, -6.975975e-13, 
    4.401784e-13, 1.345868e-13, 7.933654e-13, -2.109424e-15, -5.21444e-13, 
    -5.379724e-14, -2.825795e-12, -5.047462e-12, -3.160583e-12, -7.42395e-13, 
    -1.064371e-12, -6.383782e-13, -7.558953e-13, 3.668121e-12, 9.649448e-12, 
    5.948186e-12, 2.170153e-12, -1.664946e-12, 4.840572e-13, -9.631185e-14, 
    -2.561906e-12, -8.398837e-14, -8.973447e-13, -2.492034e-13, 
    -1.662744e-12, 1.366685e-13, 1.639577e-12, 4.004713e-14, 2.985667e-13, 
    1.654232e-13, 1.455225e-12, -4.10344e-12, -2.33763e-12, -2.387535e-13, 
    -5.278208e-13, -1.038364e-12, -6.106227e-14, 1.003642e-13, -1.337402e-13, 
    -1.49688e-12, 1.417311e-12, -2.015843e-12, -3.552825e-13, 2.443601e-13, 
    1.635797e-11, -3.762879e-13, 6.775136e-13, -2.536676e-12, 1.369401e-12, 
    -1.910812e-12, 2.203238e-13, -6.616929e-14, -3.093081e-13, -1.364631e-12, 
    -1.995404e-12, -1.125378e-12, -6.196155e-13, -6.886713e-13, 3.189116e-13, 
    1.043332e-12, 1.478706e-12, 3.718981e-12, 7.332059e-12, -2.003281e-12, 
    2.384933e-13, -3.277323e-12,
  -4.191647e-13, -1.055933e-12, 4.507505e-14, 2.498002e-15, -1.321165e-14, 
    8.277268e-13, -2.16771e-12, -2.509271e-12, -8.515744e-12, -3.121392e-13, 
    1.30479e-12, 8.312795e-13, 3.174794e-12, -4.119483e-13, 4.094614e-12, 
    -6.23307e-13, 2.577938e-13, -1.441791e-12, -1.869824e-12, -8.558154e-13, 
    -1.721567e-12, -1.220302e-12, -1.610934e-13, 1.832978e-12, -2.995382e-13, 
    -3.573419e-12, -2.294442e-12, 4.921341e-12, 2.380152e-12, -9.008128e-12, 
    -1.148748e-12, 1.929568e-13, -1.746103e-12, 3.530232e-12, -3.603562e-12, 
    -4.178213e-12, -5.400625e-13, -4.670292e-13, -2.376876e-12, 
    -9.379109e-13, -1.49436e-14, -5.848211e-12, 1.40056e-12, 6.122628e-13, 
    6.235734e-12, 5.364875e-12, -2.574052e-13, 7.684825e-13, -7.766121e-13, 
    9.352848e-12, 1.7428e-12, -2.498834e-12, 1.670591e-12, 6.115231e-12, 
    3.288245e-13, 3.805012e-13, -5.185685e-12, 3.26017e-14, -7.322032e-13, 
    1.818011e-12, -9.418466e-12, -8.301582e-12, -7.277068e-12, -8.112844e-13, 
    4.18876e-13, -2.3479e-12, 2.103595e-12, -2.625566e-12, 1.157408e-13, 
    5.75795e-12, 8.101741e-12, -5.645873e-12, 3.10274e-12, -4.23328e-13, 
    -5.450418e-12, -4.95548e-13, -6.876583e-13, -1.030495e-12, -7.978071e-12, 
    -1.307449e-11, 4.46404e-12, -1.546228e-12, 1.899231e-12, 9.638401e-13, 
    2.705169e-12, -1.123845e-11, 3.391731e-13, -8.563705e-13, -7.004597e-13, 
    -1.023015e-12, -4.42929e-12, -6.410205e-13, -1.880579e-13, -2.027884e-12, 
    -9.686696e-14, 2.062961e-12, 1.619416e-12, -3.877454e-13, 1.063355e-11, 
    4.557177e-12, -1.409428e-12, -1.524746e-12, 2.159557e-13, -2.156605e-12, 
    1.787293e-12, 1.205092e-12, -1.106892e-13, 3.185785e-13, -7.066014e-13, 
    -2.005729e-12, -1.754152e-13, 2.117195e-12, 5.385692e-13, 3.711476e-13, 
    1.738387e-12, 5.035922e-12, 1.747678e-12, 1.260488e-12, 3.041317e-13, 
    -8.960832e-12,
  -3.894329e-12, 3.71092e-13, 9.018564e-12, 5.118961e-12, 2.276901e-12, 
    -1.875333e-12, 1.152411e-13, -7.467471e-12, 1.775091e-11, 2.230127e-11, 
    -1.584677e-12, -1.367489e-11, -1.069106e-11, -8.764267e-12, 1.372119e-11, 
    2.064327e-12, -4.34347e-13, -3.646583e-12, 2.1812e-12, 1.948997e-13, 
    -1.789235e-12, -1.355693e-12, -8.980039e-13, 2.475187e-12, 4.508116e-12, 
    1.667344e-11, 1.574491e-11, 6.542489e-12, 9.484968e-12, 1.133094e-12, 
    2.177258e-12, -7.071288e-12, 1.864953e-12, 3.670064e-12, -2.253753e-14, 
    -1.657396e-12, -3.662421e-12, -6.473364e-13, -2.045392e-11, 
    -6.660561e-13, 4.613054e-12, -9.099443e-12, 1.40235e-13, -1.001491e-13, 
    1.14494e-11, 4.848955e-12, -1.369738e-13, 1.611211e-13, 3.569922e-13, 
    5.12632e-12, 7.861767e-14, -5.754952e-12, -8.03746e-14, 8.153311e-12, 
    4.349604e-13, 8.309187e-13, -1.202677e-11, 6.540102e-13, -6.305512e-13, 
    1.638989e-11, -4.851153e-11, -4.978795e-13, -8.503698e-12, -2.461476e-13, 
    -2.989409e-12, 2.267914e-11, 1.438266e-11, -1.413925e-12, 1.70407e-11, 
    2.359224e-14, -1.071976e-12, -6.432133e-12, 5.946521e-12, -4.922174e-13, 
    -8.482659e-13, -3.315126e-13, -4.985734e-13, 2.278872e-13, -1.504741e-11, 
    -2.188588e-11, 4.087536e-12, -9.35359e-12, 2.152306e-12, 1.431116e-11, 
    2.114975e-14, -5.83511e-12, 3.631262e-12, 2.443545e-12, -6.620659e-13, 
    -1.449951e-13, -1.251332e-12, -1.738936e-11, 4.49682e-13, -1.250716e-12, 
    2.011891e-12, -2.07096e-12, 1.103961e-12, 6.816325e-12, -9.55569e-13, 
    4.838064e-12, 3.847422e-12, 2.503484e-13, -4.162642e-13, -1.600213e-11, 
    1.938782e-12, 9.492407e-15, 5.535572e-13, 1.253164e-12, -3.086975e-13, 
    -3.584355e-13, 4.343526e-12, 2.265688e-12, -2.019107e-12, 1.761813e-12, 
    -1.058176e-11, 2.663403e-12, 9.184181e-13, -2.480302e-12, 8.080342e-15, 
    -2.982448e-12,
  2.892686e-12, -1.41992e-12, 1.283201e-11, 1.063749e-11, 8.51319e-13, 
    -1.070538e-11, 2.131229e-11, 3.6044e-11, 1.451744e-11, 1.394163e-11, 
    8.39312e-12, -2.632616e-12, 1.266987e-12, -3.880896e-12, -8.260059e-14, 
    2.020772e-12, -8.190498e-12, 7.54119e-13, 4.591674e-13, -1.967759e-12, 
    -5.776157e-12, -2.432055e-12, 7.28767e-12, 9.943601e-12, 1.729633e-11, 
    3.720629e-11, 1.108519e-11, -2.035894e-11, 9.51772e-12, 3.465006e-13, 
    -8.224588e-12, -4.597378e-12, 2.271683e-12, -6.53072e-12, -1.356826e-11, 
    2.275069e-12, 9.793277e-13, -9.852397e-13, 7.733708e-11, 3.987921e-13, 
    -6.014633e-13, -7.050693e-12, 3.99962e-12, 7.599534e-12, 1.318351e-11, 
    -7.803036e-12, -2.608191e-13, -8.860135e-13, -4.473866e-12, 1.819971e-12, 
    -5.848655e-13, 4.672818e-12, -2.323231e-12, 5.167866e-13, -3.106354e-12, 
    3.869405e-13, 3.654244e-12, 1.205391e-12, -2.09236e-12, 4.041628e-12, 
    -4.559408e-11, 2.248202e-12, 2.100931e-12, -4.842915e-12, -5.324819e-12, 
    3.535505e-13, -1.717571e-12, 1.225037e-11, 5.55746e-11, -3.170303e-11, 
    -9.243717e-13, 8.793521e-13, -2.376987e-13, 6.004641e-13, 7.453538e-13, 
    -6.505907e-14, -3.697528e-13, 2.300188e-12, -1.626322e-11, -6.972201e-14, 
    -5.987072e-12, 1.699458e-11, 7.486789e-13, 9.959866e-12, -7.238488e-12, 
    1.170619e-12, 6.368905e-12, 2.029155e-12, 7.306569e-14, -1.703415e-12, 
    -7.639389e-12, -3.494272e-12, 4.170692e-13, 8.927359e-13, -1.711686e-12, 
    1.084233e-12, -1.618938e-12, -5.558831e-12, -8.012369e-12, 2.781164e-12, 
    -8.4871e-13, -1.382092e-12, 4.400473e-13, -2.724217e-11, -2.704226e-12, 
    7.892575e-13, 6.533829e-12, 2.999767e-12, 2.450817e-13, -8.472667e-13, 
    -8.303358e-13, -2.626344e-12, 2.053108e-11, 8.53051e-12, -2.486594e-11, 
    -1.32086e-12, 9.132972e-14, -2.217631e-12, -2.757204e-13, 1.03817e-11,
  -8.519851e-13, 3.210543e-12, 6.152467e-12, 4.551304e-12, 1.746209e-11, 
    6.129752e-11, 3.50337e-11, 4.949208e-12, 5.542139e-11, -1.007328e-11, 
    -4.124701e-12, 3.774425e-12, -3.801331e-11, -1.298528e-11, -2.152167e-13, 
    8.380741e-13, -9.889112e-12, -2.527645e-12, 3.75075e-12, 4.16861e-12, 
    1.215361e-12, -1.455669e-12, 1.061484e-11, 2.423156e-11, -3.690098e-11, 
    -3.575751e-11, -6.339851e-11, -4.486467e-12, -8.570589e-12, 4.046358e-11, 
    2.546657e-11, 9.289847e-12, -1.058875e-12, 2.155776e-11, -2.857031e-11, 
    2.671746e-11, 1.466866e-12, -9.448831e-13, 7.557538e-11, 1.244671e-12, 
    6.179934e-12, 3.022027e-12, 6.716433e-12, 4.960686e-12, 4.631573e-12, 
    -1.625194e-11, -2.614298e-13, -4.583306e-12, -8.100498e-12, 1.978282e-12, 
    -3.353567e-13, -6.585454e-12, -1.913031e-12, 2.460143e-13, -4.876415e-12, 
    2.604306e-13, 3.823108e-12, 7.053524e-13, -5.857259e-13, -1.26585e-11, 
    -1.07061e-11, -2.903788e-13, 9.937051e-13, -5.699985e-12, -4.03636e-12, 
    -1.817491e-12, 4.20407e-11, -2.163769e-12, 1.71968e-12, 9.245216e-11, 
    9.849399e-12, -2.099459e-11, -1.434075e-11, 2.275902e-12, -9.082956e-13, 
    6.733503e-14, -2.855494e-13, -2.210916e-11, -6.951566e-12, -4.203304e-13, 
    -7.756351e-12, 2.624714e-11, -1.323802e-12, -4.662853e-11, 4.312384e-12, 
    1.064338e-11, -7.666534e-12, 1.632799e-11, -6.005621e-13, -4.436868e-12, 
    -1.649758e-11, -2.495093e-12, 1.619122e-13, -1.59715e-12, -1.037848e-11, 
    -2.189032e-12, -7.012868e-12, -1.656697e-11, -2.132594e-11, 
    -6.485368e-13, -1.607703e-11, -1.134409e-11, 1.604966e-13, -2.353861e-11, 
    -9.844348e-13, 8.318901e-13, 2.7367e-12, -2.773892e-13, -1.478817e-12, 
    -6.668055e-12, -3.672729e-12, 3.41599e-12, 1.594469e-11, 9.088674e-12, 
    -7.520207e-12, -7.505719e-13, -3.021888e-14, -2.419542e-12, 2.202554e-12, 
    6.019685e-12,
  4.767742e-12, -1.872003e-12, 4.336237e-11, 1.625433e-11, 6.513229e-11, 
    -9.297563e-13, -1.083073e-11, 5.488499e-12, -5.627887e-12, -1.100364e-11, 
    -2.220552e-11, 1.606854e-11, -8.634982e-12, -2.612155e-11, 4.221179e-12, 
    -1.206169e-12, -5.214002e-12, -5.285772e-13, 5.562238e-12, 8.196333e-12, 
    6.468548e-12, -5.723699e-12, 1.288802e-11, 1.445288e-12, -7.541245e-12, 
    -5.331391e-11, -2.433248e-11, -3.211648e-11, -2.514988e-12, 3.531686e-11, 
    1.695644e-11, 4.652045e-11, 5.086598e-12, 3.911665e-11, -1.90809e-11, 
    1.770678e-11, -1.23363e-12, -5.480338e-13, 1.84831e-11, 4.142242e-14, 
    -3.205736e-12, -2.830958e-12, 7.286588e-12, 3.314016e-14, -2.587447e-11, 
    3.073392e-11, -2.05197e-13, -6.5499e-12, 6.485923e-14, 1.270446e-12, 
    4.853284e-12, -3.00423e-11, -7.124301e-14, 7.538303e-13, -2.453966e-12, 
    4.077849e-13, 1.673606e-11, 9.217849e-13, 1.011663e-12, 7.095394e-12, 
    5.470957e-12, -5.684897e-13, -1.671829e-12, -4.795964e-12, -6.693801e-12, 
    1.042888e-12, 7.797329e-11, -1.318456e-11, -5.721279e-11, 1.638417e-10, 
    -7.830681e-12, 1.887424e-11, -3.481238e-11, 2.189499e-11, -4.978556e-12, 
    5.545564e-14, -1.622452e-13, -4.587018e-11, 8.146331e-13, 5.7504e-13, 
    -8.260337e-12, 8.005318e-12, -1.390832e-12, -3.339579e-11, 1.404321e-12, 
    -1.428652e-11, 5.7091e-12, 2.190575e-11, -3.10646e-12, -2.452205e-13, 
    -2.789685e-11, -2.960743e-12, 1.127667e-12, -2.28035e-11, -6.241785e-12, 
    4.928502e-13, -2.932932e-12, -3.835976e-11, -1.365347e-11, -4.02034e-12, 
    -6.459999e-12, -1.336154e-11, -9.111809e-13, -7.69259e-12, 8.142154e-12, 
    -4.454104e-12, -3.345546e-12, -9.647116e-12, -1.685813e-11, 
    -1.676115e-11, -1.307343e-11, 4.492184e-12, 2.817629e-11, 4.797224e-11, 
    1.080874e-11, -3.277323e-13, -1.01516e-13, -1.733601e-12, 7.187046e-12, 
    -4.344747e-12,
  1.091782e-11, 3.044387e-11, 4.432776e-11, 9.821255e-12, -1.178235e-11, 
    -4.867884e-12, -1.64464e-11, -9.435286e-11, -1.790567e-10, -4.581335e-11, 
    -4.600242e-11, 8.065826e-11, -1.047218e-11, -2.552292e-12, -3.143918e-11, 
    -2.083345e-12, -3.576173e-12, -5.180134e-12, 2.457409e-12, 1.62832e-11, 
    6.885492e-12, -1.240674e-11, 1.549583e-11, 1.378397e-11, -4.128187e-11, 
    -1.501285e-10, -3.249168e-11, -1.217249e-11, -1.275269e-11, 
    -1.867795e-11, -2.378153e-11, 4.018241e-11, 5.018508e-11, 1.295108e-11, 
    -5.700773e-11, 4.884204e-12, -1.202693e-12, -2.862433e-13, 1.242106e-11, 
    -2.403078e-12, -7.413292e-12, -1.952405e-11, 1.276554e-11, -6.366782e-13, 
    1.149081e-11, 5.617584e-11, -7.740475e-13, 1.29563e-13, 2.204193e-12, 
    7.093631e-14, 3.060149e-12, 1.108635e-11, 3.307021e-13, 5.965228e-13, 
    -4.09775e-13, 1.982303e-13, 1.000443e-10, 1.461142e-12, -5.497048e-13, 
    2.297787e-11, 6.931122e-12, -1.507305e-11, -4.845457e-12, -3.596301e-12, 
    -5.396239e-12, -3.216538e-12, 1.661941e-10, -8.648304e-12, -2.756728e-11, 
    2.271294e-12, 4.651146e-11, 9.649859e-11, 2.873468e-11, -1.797451e-13, 
    -4.368506e-12, -2.117195e-13, 6.528111e-14, -7.065598e-12, 7.253864e-13, 
    -2.183698e-12, -1.054229e-11, -1.031306e-12, 1.174949e-12, -4.628842e-11, 
    1.33793e-12, -1.255798e-10, -1.445009e-10, 2.291445e-11, -1.976679e-12, 
    4.515499e-12, -2.911893e-12, -2.031264e-13, 2.241651e-12, -7.084044e-12, 
    3.754774e-13, 1.779532e-12, -3.297895e-12, 4.827805e-12, -1.662814e-11, 
    -3.705347e-12, 2.177813e-11, 7.895046e-12, -1.892285e-12, 3.227349e-13, 
    2.95286e-11, -3.659961e-12, -6.540102e-12, -2.997591e-11, -2.874012e-11, 
    -2.77085e-11, -2.337963e-11, -4.464651e-12, 4.209089e-11, 6.235679e-11, 
    2.151945e-11, 2.396972e-13, 1.609823e-14, -3.478086e-13, 4.485828e-12, 
    -2.431844e-11,
  8.756085e-11, -6.355139e-12, -1.32967e-11, -2.631184e-11, -1.583311e-11, 
    -8.528733e-13, -4.068057e-11, -1.138258e-10, 3.907674e-11, -2.061571e-10, 
    -1.728884e-11, 4.656298e-11, -1.222871e-10, -4.650724e-12, 1.650102e-11, 
    -2.563705e-12, -6.535372e-12, -7.17415e-12, 2.26259e-11, 1.693135e-11, 
    1.821432e-12, -1.787548e-11, 4.402856e-11, 1.748424e-11, 2.561062e-11, 
    -2.673113e-10, -3.454326e-11, -3.453926e-11, -1.102229e-11, 9.830581e-12, 
    -4.902323e-11, 3.218936e-11, 1.044589e-10, -2.714029e-11, -1.565179e-10, 
    5.727485e-11, -9.18221e-13, -8.55982e-14, -3.306879e-10, -1.537859e-12, 
    -5.383072e-12, -8.586465e-12, 8.781031e-12, 3.472743e-13, 8.553536e-11, 
    6.912693e-12, 1.648126e-12, 3.610612e-12, 2.599121e-12, -2.342571e-14, 
    -8.793521e-13, 2.761369e-11, 1.687761e-13, 1.121769e-13, 3.24063e-13, 
    -4.473089e-13, 4.169953e-11, 1.306577e-12, 1.938671e-12, 1.388697e-11, 
    6.057377e-13, -4.75977e-11, 7.468248e-12, -5.723155e-12, -7.289547e-12, 
    -1.610667e-11, 1.267579e-10, 1.516764e-11, 7.933654e-12, -7.175482e-11, 
    3.958256e-11, 6.274448e-11, -5.121237e-11, -1.610867e-11, 4.578449e-12, 
    5.062617e-14, 6.325496e-14, -5.10092e-12, 2.914891e-13, -2.984146e-11, 
    -1.326872e-11, -2.910094e-12, -5.192513e-13, -2.518874e-11, 
    -1.254352e-11, 1.757827e-10, 7.957657e-11, 2.209832e-11, 8.225989e-13, 
    5.249134e-13, -1.898082e-11, -1.959366e-12, 1.815326e-12, 2.066303e-12, 
    -4.737544e-12, 9.839684e-13, -6.644774e-12, 7.8066e-11, -7.406298e-12, 
    -1.756018e-12, 6.102319e-11, 3.774199e-11, -2.402328e-12, 7.960577e-13, 
    5.645795e-11, 5.595235e-11, -2.56557e-11, -4.507927e-11, -2.621148e-11, 
    -3.540412e-11, -4.039613e-11, -1.546496e-11, 3.579892e-11, 5.222711e-11, 
    1.920109e-11, -2.442491e-14, 3.518574e-13, 4.860279e-13, 1.20276e-12, 
    -3.395506e-11,
  9.500778e-11, -4.124101e-11, -2.494649e-11, -1.968892e-11, -7.857492e-12, 
    -2.444689e-11, -5.206968e-11, -2.381533e-10, 2.153167e-12, -6.710832e-11, 
    -3.136846e-11, 1.965472e-11, -5.401815e-10, 6.552536e-13, 6.921796e-12, 
    -3.351941e-12, -8.659873e-12, -1.468603e-12, 2.535255e-11, 1.784017e-11, 
    1.147971e-13, -3.586687e-12, 6.400858e-11, -3.684097e-11, 1.051126e-10, 
    -1.233025e-10, -5.999934e-11, -4.262524e-11, -6.729262e-11, 9.701129e-13, 
    -5.992162e-11, -1.821492e-10, 1.766363e-10, -2.868594e-12, -2.847658e-10, 
    -6.092216e-11, -2.901768e-12, -5.551115e-14, -1.369218e-10, 1.512257e-12, 
    4.039924e-12, 1.950373e-11, 1.359302e-11, 5.98889e-13, 1.853497e-10, 
    -4.529155e-11, 7.130962e-12, -4.77729e-13, 2.199707e-12, -6.619705e-14, 
    7.653322e-13, 2.641909e-11, 1.343459e-12, 1.353273e-12, 3.584688e-13, 
    -7.800427e-13, -3.670819e-11, 1.18443e-12, 8.637847e-12, -1.282013e-11, 
    -2.058131e-12, -2.631251e-11, 9.592549e-12, -5.505951e-12, -5.396527e-12, 
    1.314755e-10, 1.672935e-10, 1.093035e-10, 1.029095e-10, 2.496292e-11, 
    2.569478e-11, 9.906809e-11, -2.793719e-10, 3.888001e-13, 1.412603e-11, 
    8.26228e-13, -1.165734e-15, -5.356049e-12, -1.45437e-12, -1.446865e-11, 
    -1.394573e-11, 1.974976e-12, -3.150813e-12, -5.618239e-11, -1.162948e-10, 
    1.702725e-10, 1.205718e-10, 2.511436e-11, 8.59382e-14, -8.553158e-13, 
    -1.268341e-11, 4.11684e-12, 8.280043e-13, -1.838991e-11, -1.982037e-11, 
    -2.805134e-12, -1.044271e-11, 3.278999e-11, 1.019185e-13, -9.984458e-13, 
    1.032705e-10, 7.09513e-12, -1.819656e-12, 1.10853e-12, 6.86462e-11, 
    1.450282e-10, -9.721401e-11, -1.210598e-10, -3.532397e-11, -2.955169e-11, 
    -4.345346e-11, -2.01672e-11, 2.237566e-11, 1.053535e-11, 1.463873e-11, 
    -1.653344e-13, 9.456325e-13, 1.659645e-13, -8.493206e-14, -1.394305e-10,
  2.45346e-11, -3.322365e-11, 1.137712e-11, -4.025624e-11, -6.203349e-11, 
    -5.174039e-11, -4.771694e-11, -3.124465e-10, -8.443868e-11, 7.07745e-12, 
    -1.307758e-10, 7.654632e-11, -6.247665e-10, 7.296386e-13, 3.996803e-15, 
    -2.907452e-12, -8.443734e-12, 1.018652e-11, 2.144662e-11, 2.832001e-11, 
    -4.60032e-12, 2.291722e-11, 4.323431e-11, -9.936807e-11, -6.283418e-12, 
    1.011524e-10, -1.057567e-10, -5.137002e-11, -1.655365e-10, -4.606315e-11, 
    -8.118528e-11, -6.406031e-11, 1.818123e-10, -3.301581e-11, -5.073053e-11, 
    -1.881966e-10, -6.868816e-12, -1.898481e-13, 3.950764e-10, 5.197442e-12, 
    5.806466e-12, 4.045697e-11, 3.813194e-11, -2.712677e-12, -1.804898e-10, 
    -2.262204e-10, 1.827827e-11, 1.275957e-11, 2.18483e-12, -4.591882e-13, 
    -3.324563e-12, 3.894618e-11, 7.891643e-12, 5.854072e-12, -1.939782e-13, 
    2.398082e-14, -3.70854e-10, 2.006484e-12, 1.566907e-11, -5.718537e-11, 
    3.429701e-12, 9.866641e-11, 1.89071e-11, 3.693934e-13, 4.459811e-12, 
    1.080962e-10, 2.989773e-10, 2.599143e-10, 1.230336e-10, 1.194747e-10, 
    -2.828626e-11, 4.675162e-10, 2.817715e-10, 8.194911e-11, 1.70556e-11, 
    2.07967e-12, 1.068035e-13, -3.23408e-12, -3.564615e-12, 1.045071e-10, 
    -1.356115e-11, 7.668954e-12, -6.12177e-12, -5.959189e-11, -9.044454e-11, 
    -2.895351e-10, -1.636811e-10, 3.088596e-11, -3.008302e-12, 3.173906e-12, 
    -4.586598e-11, -1.790648e-11, 4.143352e-13, -3.489671e-11, -5.46474e-11, 
    -1.354321e-11, -1.752243e-11, 2.505418e-11, 3.006484e-13, 2.675637e-12, 
    1.239671e-10, 1.986189e-10, -8.334444e-13, 1.14958e-12, 2.293588e-11, 
    1.929927e-10, -7.709255e-11, -2.596106e-10, -5.636869e-11, -2.263301e-11, 
    -3.869305e-11, -1.26632e-11, -2.48912e-12, -2.710854e-11, 1.124745e-11, 
    -1.713296e-13, 1.763034e-12, -2.96041e-13, -7.875367e-13, -1.110423e-10,
  -1.836309e-12, 1.402878e-12, 2.108669e-11, -7.35545e-12, -5.80731e-11, 
    -2.274314e-11, -7.352563e-11, -2.995333e-10, -3.38011e-10, -1.425717e-10, 
    -8.175371e-11, 2.658846e-10, -9.475269e-10, 2.577716e-11, -2.823652e-11, 
    -8.458123e-13, -3.939959e-12, 1.753664e-11, 3.651934e-11, 3.673994e-11, 
    -1.42939e-11, 2.273248e-11, -1.961764e-11, -2.068048e-10, 3.944356e-11, 
    -9.648149e-11, -1.669114e-10, -4.735279e-11, -3.790244e-10, 
    -4.640599e-11, -2.305129e-10, -4.992406e-11, 2.016285e-10, -2.155516e-10, 
    2.36748e-10, -4.53714e-10, -1.153939e-11, -2.853273e-13, 8.55239e-10, 
    2.14647e-11, -8.150449e-11, 3.422818e-11, 6.375567e-11, -1.135149e-11, 
    3.555822e-12, -5.760925e-10, 3.518652e-11, 9.177126e-11, 4.697576e-13, 
    -1.10556e-12, 1.511369e-11, 1.125167e-10, 2.333858e-11, 2.833378e-12, 
    -2.743139e-13, -6.794565e-14, 7.173049e-10, 2.212808e-12, 2.673204e-11, 
    -9.729129e-11, 1.023226e-11, 1.727645e-10, -1.820366e-11, 9.778756e-12, 
    1.435678e-11, 1.291247e-10, 6.156986e-11, 4.044876e-10, 2.134972e-10, 
    1.840497e-10, -1.163136e-10, 8.713665e-10, 2.514846e-10, 1.3141e-10, 
    1.7174e-11, 2.291944e-12, 2.14051e-13, 2.705836e-12, -1.872547e-12, 
    2.418497e-10, -1.709033e-11, 1.011147e-11, -9.844126e-12, -1.562062e-10, 
    -8.951551e-11, -1.056646e-09, -1.071809e-11, 3.701706e-11, -8.963844e-12, 
    1.063016e-11, 7.080425e-11, -4.862182e-11, 6.705747e-13, -3.14035e-11, 
    -6.89675e-11, -3.089031e-11, -3.356506e-11, 1.993516e-12, -4.264589e-12, 
    6.406342e-12, 2.401239e-10, 6.454852e-10, 2.426948e-13, 2.428835e-12, 
    -1.825651e-12, 7.968159e-11, 1.248295e-10, -3.0369e-10, -5.046763e-11, 
    -1.230527e-11, -2.721423e-11, 5.990763e-13, -3.342526e-11, -7.832446e-11, 
    1.326894e-11, -1.528555e-13, 2.695622e-12, -3.799183e-13, -2.29472e-12, 
    1.298672e-10,
  -2.865796e-11, 3.146461e-11, 1.858158e-10, 2.213696e-10, 7.398704e-11, 
    -4.866507e-11, -1.679794e-10, -2.721237e-10, -5.184884e-10, -7.65823e-11, 
    4.679617e-10, 1.149102e-09, -8.470504e-10, 7.055334e-11, -2.48388e-11, 
    3.844747e-12, 4.508216e-12, 1.579537e-11, 6.92264e-11, 3.104006e-11, 
    -2.71676e-11, 1.820766e-11, -9.512924e-11, -3.023803e-10, 1.889937e-10, 
    -5.758167e-10, -1.587921e-10, 1.133866e-10, -7.997087e-10, -8.386181e-11, 
    -2.305143e-10, 4.410161e-11, 1.721823e-10, -9.785417e-11, 4.342233e-10, 
    -7.553815e-10, -1.424265e-11, -5.906386e-14, 1.54326e-09, 8.141647e-11, 
    -2.059405e-10, 6.949108e-12, 6.42566e-11, -1.960418e-11, 3.490577e-10, 
    -9.430714e-10, 5.573142e-11, 2.219451e-10, -9.005419e-12, -1.798561e-12, 
    3.775025e-11, 3.560494e-10, 4.756746e-11, -2.049596e-11, 3.707612e-12, 
    -4.316547e-13, 2.432968e-09, 4.311573e-12, 3.625882e-11, -5.031864e-11, 
    2.0421e-11, 1.709175e-10, 6.981082e-13, 1.43519e-11, 1.681748e-11, 
    2.183853e-11, -1.058318e-10, 1.650236e-10, 3.936851e-10, 2.347562e-10, 
    -1.049756e-10, 1.91808e-09, 2.098872e-10, 1.519069e-10, 1.26068e-12, 
    -2.611245e-13, 2.664535e-13, 1.483746e-11, 5.215961e-12, 4.036735e-10, 
    -3.559553e-11, 1.203069e-11, -1.016698e-11, -2.152429e-10, -8.425793e-11, 
    -1.870232e-09, 1.651905e-10, 4.444978e-11, -2.455619e-11, -1.054978e-11, 
    4.279599e-10, -2.704077e-11, -2.651213e-13, -2.624514e-11, -3.737455e-11, 
    -5.557936e-11, -5.574101e-11, 2.17959e-11, -1.142375e-11, 7.753442e-12, 
    5.868515e-10, 8.970802e-10, 1.923128e-12, 9.487966e-12, 7.714362e-11, 
    1.271392e-10, 3.367777e-10, -3.477307e-10, -8.846968e-11, -7.716494e-12, 
    -1.094413e-11, 8.526513e-12, -6.159873e-11, -1.239115e-10, 1.520561e-11, 
    6.181722e-13, 2.712497e-12, -8.187895e-14, -4.910405e-12, 3.083294e-10,
  -5.317702e-11, -5.041656e-11, 7.50191e-11, 3.535519e-10, 5.410925e-10, 
    2.02359e-10, -3.990728e-10, -3.402576e-10, -2.857341e-10, 8.580905e-10, 
    1.491241e-09, -3.602345e-10, -5.845173e-10, 1.208669e-10, 4.436274e-11, 
    1.004388e-11, 1.646825e-11, 1.209344e-11, 1.026246e-10, 1.719869e-11, 
    -3.530332e-11, 3.502265e-11, -1.188667e-10, -2.189431e-10, 4.558274e-10, 
    3.380016e-10, -3.324097e-10, 4.41112e-10, -1.834316e-09, -2.338716e-10, 
    -6.110525e-10, 1.420872e-10, 1.075229e-10, -9.783534e-10, 2.334346e-10, 
    -8.576926e-10, -2.528466e-11, 1.414424e-12, 4.205233e-09, 2.142897e-10, 
    5.703314e-11, -5.267609e-11, 5.281642e-11, -2.208839e-11, 1.923617e-10, 
    -1.059988e-09, 8.22169e-11, 2.411058e-10, -2.474678e-11, -4.575895e-12, 
    -4.265566e-11, 1.086104e-09, 9.974279e-11, -4.15632e-11, 1.156204e-11, 
    -1.172396e-12, 3.891319e-09, 1.563976e-11, 5.122622e-11, 1.654885e-10, 
    1.242029e-11, 1.332161e-10, -3.267786e-11, 1.751346e-11, 1.402398e-11, 
    9.385204e-11, -1.646328e-09, -2.579768e-10, 6.416521e-10, 2.613234e-10, 
    1.317595e-10, 4.403098e-09, -2.476632e-10, 2.361595e-10, 2.722196e-11, 
    -2.973621e-12, 6.261658e-13, 3.190959e-11, 1.016742e-11, 5.66807e-10, 
    -9.131718e-11, 1.58602e-11, -2.881251e-12, -3.005063e-10, -6.548007e-11, 
    -1.922444e-09, -7.194245e-12, 4.616396e-11, -6.700218e-11, -1.186571e-10, 
    8.016805e-10, 8.671677e-11, -3.662848e-12, -9.083934e-12, -1.851603e-10, 
    -7.92447e-11, -7.544472e-11, 2.058869e-10, -2.22613e-11, 6.554046e-12, 
    9.148273e-10, 7.9621e-10, 4.414469e-12, 2.732858e-11, 1.162626e-10, 
    2.440146e-10, 3.008651e-10, -7.539249e-10, -6.484235e-10, -2.861e-11, 
    5.428547e-12, -1.184475e-11, -1.041762e-10, -2.067964e-10, 2.502887e-11, 
    2.478018e-12, 2.470912e-12, 4.458656e-13, -5.550671e-12, 3.078107e-10,
  1.426059e-11, 2.300382e-11, -4.43876e-11, -5.240963e-11, 5.211724e-10, 
    8.101786e-10, -2.144951e-10, -5.160778e-10, -1.940883e-10, 2.547296e-10, 
    8.871659e-10, 5.211476e-11, 4.509957e-10, 1.934346e-10, 1.973142e-10, 
    8.654411e-12, 2.815028e-11, 1.184119e-11, 1.217222e-10, 1.408296e-11, 
    -3.478107e-11, 6.0421e-11, -1.237339e-10, -1.610978e-10, 1.38008e-09, 
    1.841837e-09, -7.970016e-10, -5.190088e-10, -2.213152e-09, -7.02876e-10, 
    -1.475321e-09, 2.479688e-10, -4.788667e-10, -1.391779e-09, 6.33591e-11, 
    -1.383121e-09, -3.976197e-11, 4.439116e-12, 5.940034e-09, 3.552817e-10, 
    3.579622e-10, -1.453415e-10, 4.507417e-11, -2.212031e-11, 4.42153e-10, 
    -9.443433e-10, 1.33344e-10, -2.825118e-11, -3.858602e-11, -1.232103e-11, 
    -1.942868e-10, 1.280213e-09, 2.777213e-10, -5.598935e-11, 1.698037e-11, 
    -2.31104e-12, 6.062042e-09, 3.601883e-11, 1.697252e-10, 3.035683e-10, 
    -4.973799e-12, 7.18039e-11, 9.604051e-11, 2.36362e-11, 1.56092e-11, 
    8.93813e-10, -9.66633e-10, -5.631193e-10, 9.059917e-10, 2.659384e-10, 
    3.406839e-10, 5.196306e-09, 7.357528e-10, 3.875655e-11, 5.209344e-11, 
    -1.275424e-12, 1.642242e-12, 3.92788e-11, 1.328333e-11, 7.783889e-10, 
    -1.722498e-10, -5.614104e-11, 4.382272e-12, -3.313261e-11, 7.460699e-12, 
    7.369287e-10, -5.433733e-10, 6.149037e-11, -1.725065e-10, -1.930864e-10, 
    6.675194e-10, 3.929436e-10, -7.72804e-12, -3.709388e-11, -2.548859e-10, 
    -9.350565e-11, -1.025569e-10, 5.605827e-10, -3.21414e-11, 4.455814e-12, 
    8.564633e-10, 5.987231e-10, 4.877876e-12, 5.016765e-11, -8.504131e-11, 
    2.038263e-10, -8.619949e-11, -1.131511e-09, -1.218552e-09, -1.180211e-11, 
    2.336975e-11, -5.019984e-11, -2.387104e-10, -3.377387e-10, 3.41096e-11, 
    4.781953e-12, 4.045653e-12, 9.342527e-13, -4.020118e-12, 1.950902e-10,
  2.461498e-10, 2.740315e-10, 2.803517e-10, 9.987389e-11, 1.00755e-10, 
    6.842988e-10, 5.600818e-10, -6.103242e-10, -4.867822e-10, -6.215899e-10, 
    -9.145396e-11, 9.800871e-11, 7.334151e-10, 3.580034e-10, 4.957954e-10, 
    -2.641762e-11, 2.57252e-11, 1.776179e-11, 1.174647e-10, 1.679723e-11, 
    -3.935341e-11, 4.938983e-11, -3.177973e-10, -7.397176e-10, 2.593772e-09, 
    8.924737e-10, -1.370562e-09, -2.136947e-09, -1.215675e-09, -1.680942e-09, 
    -2.537707e-09, 6.082814e-10, -7.607923e-10, -1.8651e-09, 2.25775e-11, 
    -1.559762e-09, -5.23837e-11, 8.686385e-12, 5.884914e-09, 2.891273e-10, 
    6.354881e-11, -1.801794e-10, 7.07665e-11, -2.425282e-11, 3.087628e-10, 
    -7.83043e-10, 2.376321e-10, -4.577254e-10, -4.348948e-11, -2.851208e-11, 
    -1.480469e-10, 5.307648e-10, 7.190493e-10, -7.624266e-11, 2.88896e-11, 
    -3.581135e-12, 7.368328e-09, 4.788845e-11, 6.920128e-10, 1.291975e-10, 
    -2.043521e-11, 3.730349e-12, 4.592096e-10, 2.709584e-11, 2.804583e-11, 
    7.591439e-10, 4.664713e-12, -9.541452e-10, 1.443826e-09, 9.914558e-11, 
    1.399698e-10, 5.862493e-09, -1.511253e-10, -3.979217e-10, 1.621991e-10, 
    6.82121e-12, 2.753353e-12, 6.907008e-11, 2.29555e-11, 9.580283e-10, 
    -2.143885e-10, -1.517074e-10, 1.002221e-11, -7.954242e-10, 9.27507e-11, 
    2.095472e-09, -2.811582e-10, 1.012346e-10, -3.827e-10, 1.049028e-10, 
    5.052634e-10, 8.566566e-10, -8.373746e-12, -3.808864e-11, -4.126974e-10, 
    -8.556391e-11, -1.654044e-10, 1.150724e-09, -2.666667e-11, 2.231104e-13, 
    6.370335e-10, 5.248584e-10, 1.289191e-12, 6.550893e-11, -6.259206e-10, 
    6.750511e-11, -6.503598e-11, -1.166736e-09, -4.645919e-10, 5.348504e-10, 
    6.253842e-11, -6.465228e-11, -3.896581e-10, -4.449277e-10, 3.084821e-11, 
    9.954704e-12, 1.12288e-11, 2.016165e-13, 1.736389e-13, 9.972823e-11,
  4.367031e-10, 8.286953e-10, -2.063434e-09, -1.117009e-10, 2.8108e-10, 
    1.015827e-10, 1.090367e-09, -5.57133e-10, -7.353655e-10, -7.262564e-10, 
    6.991066e-10, -6.520899e-10, 9.406129e-10, 6.082566e-10, 9.535519e-10, 
    -1.785743e-10, -1.021405e-11, 4.611422e-12, 1.101368e-10, 2.113509e-11, 
    -5.971046e-11, -1.277911e-11, -4.447749e-10, -2.09192e-09, 2.82861e-09, 
    -1.50332e-09, -9.196874e-10, -2.762651e-09, -2.168466e-09, -4.057863e-09, 
    -3.268372e-09, 4.780425e-10, -1.274838e-09, -3.77273e-09, 8.853007e-11, 
    -1.852438e-09, 2.250431e-11, 9.257484e-12, 6.275879e-09, -1.671999e-10, 
    -1.327471e-10, -7.549161e-11, 2.082441e-10, -2.514033e-11, -2.061793e-09, 
    -6.334382e-10, 3.708607e-10, -4.765539e-10, -4.191136e-11, -3.232969e-11, 
    -9.355006e-11, -1.06791e-10, 1.350873e-09, 9.872991e-12, 1.206587e-10, 
    -5.002221e-12, 2.798874e-09, 3.466951e-11, 1.954972e-09, 7.709389e-13, 
    -3.61986e-11, -7.596057e-11, 2.430092e-10, 1.001226e-11, 3.335643e-11, 
    -8.041035e-10, 2.023942e-09, -5.970939e-10, -9.903864e-10, -7.203838e-11, 
    1.16021e-10, 4.727351e-09, -2.471587e-10, -8.058159e-10, 6.755627e-10, 
    1.914557e-11, 9.672263e-13, 2.26736e-10, 5.512604e-11, 9.212364e-10, 
    -2.080967e-10, -4.295078e-10, 1.090683e-11, -1.798135e-10, 1.095977e-10, 
    1.400604e-09, 8.304077e-10, 1.482299e-10, -7.489062e-10, 5.901057e-10, 
    6.581722e-10, 1.364034e-09, -6.696865e-12, 8.903598e-11, -8.82391e-10, 
    -4.313705e-11, -2.554834e-10, 1.50548e-09, -5.318412e-12, -9.446666e-12, 
    5.375256e-12, 6.569794e-10, -1.597389e-12, 8.328138e-11, -1.222237e-09, 
    -4.741914e-10, 2.126548e-10, -1.613866e-09, -1.049436e-10, 1.395588e-09, 
    1.623199e-10, -1.286189e-10, -4.83606e-10, -5.669598e-10, 2.877343e-11, 
    1.776286e-11, 5.158629e-11, -5.730971e-12, 2.575717e-12, 1.708855e-12,
  4.540475e-10, 8.982362e-10, -3.321606e-09, -5.144617e-09, -6.075318e-10, 
    1.105786e-09, 7.035901e-10, 5.355751e-10, -8.598882e-10, 3.105605e-10, 
    2.619455e-09, -2.213969e-09, 1.259988e-09, 9.451178e-10, 1.053191e-09, 
    -5.583125e-10, -1.614516e-10, -3.812062e-12, 1.335394e-10, 4.675016e-11, 
    -1.075797e-10, -9.477574e-11, -3.86752e-10, -2.51892e-09, -5.366623e-10, 
    -4.344063e-09, 9.018883e-10, -1.384311e-09, -2.778297e-09, 1.859473e-09, 
    -5.830604e-09, 1.342894e-09, -4.54552e-10, -3.739448e-09, 3.503082e-10, 
    -3.223096e-09, 2.210548e-10, 2.680522e-12, 2.629999e-09, -5.033833e-10, 
    2.712781e-11, 1.171507e-10, 5.394689e-10, -1.266698e-10, -3.054485e-09, 
    -5.131575e-10, 5.00247e-10, 2.272316e-11, -1.110784e-10, -4.051426e-11, 
    -2.524398e-10, -1.564224e-10, 1.855387e-09, 1.727948e-10, 3.718625e-10, 
    -6.526335e-12, 5.178684e-10, 1.172609e-11, 3.757328e-09, 2.490221e-10, 
    -4.707346e-12, -2.679919e-10, 6.46132e-11, 3.756426e-11, 2.101999e-11, 
    -2.740709e-09, -5.299785e-09, 3.943622e-09, 1.314103e-09, -4.961365e-11, 
    1.862581e-10, 2.364256e-09, 6.440004e-11, -9.75394e-10, 8.758739e-10, 
    4.108003e-11, -1.8332e-12, 5.458993e-10, 8.266383e-11, -4.060396e-11, 
    -2.89166e-10, -7.547687e-10, 3.673861e-11, -1.58412e-10, 1.404281e-10, 
    -1.427516e-10, 1.657408e-09, 1.780158e-10, -1.284034e-09, 6.614407e-10, 
    9.465957e-10, 1.92563e-09, -2.973621e-12, 1.320792e-10, 1.239862e-10, 
    4.52971e-12, -3.142823e-10, 1.977977e-09, 2.240697e-11, -3.142944e-11, 
    -5.910756e-10, 8.793322e-10, -3.081979e-12, 1.161444e-10, -1.473143e-09, 
    -1.546258e-09, -1.320007e-09, -6.869421e-10, 7.15481e-11, 1.529155e-09, 
    6.310152e-10, -3.246079e-10, -6.000995e-10, -7.226539e-10, 5.679723e-11, 
    2.736371e-11, 1.343885e-10, -2.218803e-11, -5.815792e-12, -1.502265e-10,
  -5.390532e-11, 2.332197e-09, 2.788394e-09, -5.469904e-09, -5.079517e-09, 
    8.117205e-10, -1.176975e-09, 1.806679e-09, 1.006224e-09, 2.49997e-09, 
    4.301338e-09, -2.286473e-09, 1.487415e-10, 1.223167e-09, 1.796121e-09, 
    -1.002446e-09, -3.132207e-10, -2.876632e-11, 1.998846e-10, 1.491536e-10, 
    -1.810356e-10, -1.858105e-10, -2.629328e-10, -1.130292e-09, -6.46553e-09, 
    -2.549474e-09, 2.922459e-09, 7.513528e-10, -3.095526e-09, 3.362214e-09, 
    -6.985761e-09, 3.123795e-10, 1.936396e-09, -1.760331e-09, 7.365735e-10, 
    -4.77009e-09, 3.277386e-10, 8.79119e-12, 5.020066e-09, 5.840306e-11, 
    5.453636e-10, 3.086242e-11, 8.807106e-10, -4.996417e-10, -2.964331e-09, 
    -1.811067e-10, 6.515357e-10, 4.9031e-10, -5.111431e-11, -4.417178e-11, 
    -2.81716e-10, -1.174847e-10, 2.194043e-09, 2.839919e-10, 5.829947e-10, 
    -6.703971e-12, -1.621945e-09, 1.852314e-11, 5.339674e-09, -3.742144e-10, 
    6.283685e-11, -4.314025e-10, -2.592415e-11, 9.413661e-10, 7.229773e-12, 
    -4.45127e-09, -7.750717e-09, 3.008221e-09, 3.154678e-09, 1.113243e-10, 
    -2.311431e-10, 4.334918e-09, 1.903224e-10, -1.690843e-10, 2.84836e-10, 
    3.94742e-11, 7.496226e-12, 8.659171e-10, 2.807923e-11, 8.979484e-11, 
    -6.999166e-10, -2.509186e-10, 1.422968e-10, 6.959137e-09, 7.033627e-10, 
    -1.881695e-10, 1.610925e-09, 1.786553e-10, -1.868502e-09, 3.756178e-10, 
    9.90422e-10, 2.792381e-09, 1.148592e-11, 4.243859e-11, -6.601404e-10, 
    1.996838e-11, -3.404729e-10, 2.58559e-09, 6.542322e-11, -6.381029e-11, 
    -9.167316e-10, 7.998411e-10, -7.842615e-12, 1.510321e-10, -1.64032e-09, 
    -3.788532e-09, -3.932531e-09, -3.148461e-09, -1.621476e-09, 2.52933e-09, 
    1.674916e-09, -4.675407e-10, -6.232206e-10, -1.004839e-09, 6.292211e-11, 
    3.095053e-11, 2.329905e-10, -4.166756e-11, -4.991652e-11, -3.0089e-10,
  -1.109036e-09, -1.059469e-09, -3.112596e-09, -2.431896e-09, -5.881411e-09, 
    -6.179555e-09, -5.689387e-10, 1.826415e-09, 2.636092e-09, 3.692072e-09, 
    4.969202e-09, 3.425136e-09, 5.566179e-10, 1.620414e-09, 2.6536e-09, 
    -6.658767e-10, -2.764821e-10, -1.237055e-11, 2.823306e-10, 2.358789e-10, 
    -2.219664e-10, -3.275815e-10, -3.867484e-11, 2.128004e-10, -2.635254e-09, 
    5.939356e-10, 3.767653e-10, 1.692584e-10, -5.182436e-09, -6.442541e-09, 
    -8.48825e-09, -1.440689e-09, 5.058816e-09, -1.433953e-09, 9.557439e-10, 
    -5.6095e-09, -4.28173e-12, 1.901768e-11, 7.049302e-09, 3.423068e-10, 
    1.283617e-09, -4.32884e-10, 2.060631e-09, -5.812986e-10, -2.517559e-09, 
    4.347456e-10, 8.085621e-10, 9.368861e-10, 3.239805e-10, -6.988543e-11, 
    -1.908909e-10, -4.180478e-10, 2.501231e-09, 3.401809e-10, 5.748881e-10, 
    -1.090683e-11, -5.452499e-09, 7.930936e-11, 5.842479e-09, -7.309694e-09, 
    1.47601e-10, -4.560476e-10, 5.650946e-11, 4.221279e-09, -1.324899e-09, 
    -2.670781e-09, -6.559468e-09, 2.30731e-09, 6.170048e-09, 2.375558e-10, 
    -7.531966e-10, 5.3249e-09, 3.809717e-10, -7.718413e-10, 1.309458e-09, 
    3.765876e-13, 6.494361e-12, 8.384404e-10, 4.974652e-11, -1.472152e-09, 
    -1.074021e-09, 7.348375e-10, 3.58888e-10, 7.935981e-10, -2.346709e-10, 
    -5.217515e-11, 6.53479e-10, 1.665583e-10, -2.476798e-09, 3.686935e-10, 
    6.951169e-10, 4.130807e-09, 1.089262e-11, -3.257739e-10, 8.111911e-10, 
    2.330722e-11, -4.09328e-10, 2.686654e-09, 1.431957e-10, -8.117098e-11, 
    4.110419e-10, 2.666205e-10, -2.043876e-11, 1.663807e-10, -2.872746e-09, 
    -3.876089e-09, -4.55767e-09, -5.211881e-09, -2.286633e-09, 5.562903e-09, 
    3.579352e-09, -4.110845e-10, -2.966871e-10, -1.456804e-09, -7.465673e-11, 
    2.147118e-11, 2.532268e-10, -3.403322e-11, -9.083578e-11, -3.725162e-10,
  -2.876277e-09, 1.953993e-10, 1.097789e-09, -5.516341e-09, -9.403323e-09, 
    -1.288777e-08, 2.643532e-09, 6.11351e-10, 3.383093e-09, 3.921912e-09, 
    4.978887e-09, 7.033492e-09, 3.103651e-11, 1.203915e-09, 2.962764e-09, 
    -7.822964e-10, -6.946607e-10, 4.95902e-10, 5.755396e-12, 8.341772e-10, 
    -1.958824e-10, -4.847038e-10, -1.286367e-10, 1.256808e-09, 8.099079e-09, 
    2.747186e-09, -9.07346e-09, -9.387406e-10, -1.51465e-09, -2.889337e-08, 
    -1.141652e-08, -4.092669e-09, 5.311989e-09, -1.06894e-09, 5.907452e-10, 
    -8.313549e-09, -2.842284e-10, 5.94369e-12, 4.800768e-09, 9.198855e-10, 
    1.999029e-09, -9.410712e-10, 4.317613e-09, -6.808087e-10, 7.614176e-11, 
    6.902781e-10, 8.811298e-10, 1.199027e-09, 5.174399e-10, -1.381242e-10, 
    3.177192e-11, -8.105303e-10, 2.996288e-09, 4.254332e-10, 6.726715e-10, 
    -3.616663e-11, -1.220741e-09, 1.885184e-10, 2.715871e-09, -8.452904e-09, 
    2.148397e-10, -6.333494e-10, 1.606963e-10, 7.258666e-09, -3.86824e-09, 
    -1.012353e-09, -5.049827e-09, 1.37527e-09, 4.840871e-09, 7.514984e-10, 
    -1.427594e-09, 1.228238e-08, 6.890843e-10, -2.494005e-09, 2.609767e-09, 
    -1.045919e-11, -1.599787e-11, 7.692549e-10, 1.883777e-10, -4.133511e-09, 
    -1.68663e-09, 6.172023e-10, 5.447731e-10, 6.069541e-09, 5.773387e-09, 
    -7.42773e-10, 1.467669e-09, 8.489565e-11, -2.278021e-09, 3.762182e-10, 
    7.833307e-10, 5.591068e-09, 1.98952e-12, -2.51128e-09, 1.819274e-09, 
    5.11875e-11, -5.502386e-10, 1.778488e-09, 2.957563e-10, -5.689458e-11, 
    1.744752e-09, -3.81144e-10, -2.725642e-11, 2.03956e-10, -3.444768e-09, 
    -1.044981e-09, -3.250022e-09, -6.37877e-09, -3.193293e-09, 7.711407e-09, 
    6.219466e-09, -6.525909e-10, 5.704237e-11, -2.384013e-09, -2.657146e-10, 
    -1.69706e-11, 1.240963e-11, 3.181633e-11, -1.079723e-10, -4.8027e-10,
  -3.903551e-09, 2.187249e-09, 3.359588e-09, -2.881762e-09, -6.337018e-09, 
    -6.937398e-09, 1.713545e-10, -8.472512e-10, 2.876419e-09, 4.316973e-09, 
    3.523866e-09, 1.248549e-08, -3.040839e-10, -1.690466e-09, 4.307594e-10, 
    2.940115e-10, -1.039862e-09, -1.029008e-10, -4.050342e-10, 3.090918e-09, 
    -9.229382e-10, -7.404992e-10, -3.243485e-10, 5.595666e-10, 9.11848e-09, 
    5.136712e-09, -1.808326e-08, -5.057416e-09, 1.117269e-08, -3.463532e-08, 
    -1.709509e-08, -3.371099e-09, -4.093579e-10, -6.757546e-10, 
    -1.290346e-11, -1.138645e-08, -4.177309e-10, 1.190159e-12, -1.625097e-09, 
    1.602424e-09, 2.330427e-09, -1.432539e-09, 5.938965e-09, -1.106545e-09, 
    2.662745e-09, 1.197606e-09, 1.299156e-09, 1.916533e-09, 1.642218e-09, 
    -2.984404e-10, 4.455245e-10, -6.183711e-10, 3.763611e-09, 2.515606e-10, 
    1.165415e-09, -9.811174e-11, 1.61441e-09, 3.151939e-10, 1.343287e-09, 
    -9.605881e-09, -6.662049e-11, -1.153552e-09, -6.361915e-10, 8.447034e-09, 
    -1.831154e-09, 6.782074e-09, -3.910742e-09, 2.309548e-10, 7.8293e-09, 
    1.139767e-09, -2.774868e-09, 2.048688e-08, 4.375238e-10, -1.345995e-09, 
    2.801627e-09, 6.400569e-11, -7.479528e-11, 1.315875e-09, 3.282181e-10, 
    9.496262e-10, -1.67951e-09, 2.160476e-10, 5.525322e-10, 5.399556e-09, 
    5.051419e-09, -6.287735e-10, 3.135796e-09, -9.896439e-11, -1.315642e-09, 
    2.615934e-10, 3.872231e-09, 6.411972e-09, -6.445333e-11, -9.72013e-09, 
    2.587512e-09, 2.578702e-10, -5.537572e-10, 6.678533e-10, 3.639116e-10, 
    3.400373e-11, 2.494346e-09, -9.476917e-10, 4.364509e-12, 2.962803e-10, 
    -1.808985e-09, -2.413003e-11, -2.26413e-09, -3.437236e-09, -1.122913e-09, 
    8.269694e-09, 6.611941e-09, -1.245638e-09, 2.137313e-11, -3.458041e-09, 
    -3.708465e-10, -6.259597e-11, -4.49333e-10, 9.147882e-11, -1.111431e-10, 
    -5.226468e-10,
  -2.11196e-09, 1.3072e-09, 3.506074e-09, 1.569163e-09, -3.386873e-09, 
    -1.858211e-09, -1.171253e-08, -1.308138e-09, 2.070465e-09, 3.100837e-09, 
    3.268553e-09, 9.974997e-09, -2.070237e-10, 2.802864e-09, 1.459597e-09, 
    1.306271e-09, -2.197606e-09, -1.547889e-09, -4.031477e-10, 5.742692e-09, 
    -2.596522e-09, -1.347871e-09, -4.998526e-10, -4.439471e-11, 7.534595e-10, 
    1.363796e-08, -1.841804e-08, -8.346973e-09, 2.136389e-08, -1.920765e-08, 
    -2.479021e-08, -7.993606e-10, -3.786909e-09, -1.916476e-10, 
    -1.050751e-10, -1.207897e-08, -9.135789e-10, -6.465939e-11, 
    -5.347232e-09, 2.435885e-09, 2.102513e-09, -2.159368e-09, 6.882637e-09, 
    -1.921179e-09, 1.020047e-08, 2.176478e-09, 1.662215e-09, 3.432504e-09, 
    3.491567e-09, -5.23757e-10, 1.059117e-09, -1.232934e-10, 4.912391e-09, 
    -1.59713e-10, 3.820885e-09, -1.328999e-10, 2.662404e-09, 4.339711e-10, 
    -4.899334e-11, -1.338681e-08, -1.614353e-09, -1.105434e-09, 
    -1.463633e-09, 2.047392e-09, -1.3288e-09, 1.25618e-08, -2.689035e-09, 
    1.13468e-09, 1.217154e-08, -4.715162e-10, -2.726352e-09, 8.283592e-09, 
    -5.968843e-10, 5.541096e-10, 4.337639e-09, 7.810286e-11, -1.911893e-10, 
    1.457778e-09, 4.164512e-10, 9.866113e-09, -2.694051e-09, -5.519931e-10, 
    3.197442e-10, 2.585324e-09, 2.396405e-09, 1.829449e-09, 2.171873e-09, 
    -2.463025e-10, -1.901412e-11, 6.146195e-11, 8.459523e-09, 6.61874e-09, 
    -2.979377e-10, -2.634019e-08, -8.036238e-10, 7.224514e-10, -8.35314e-11, 
    1.022528e-09, 5.55417e-10, -3.268497e-11, 2.571568e-09, -1.407155e-09, 
    9.382539e-11, 4.05965e-10, -7.372307e-10, 2.621903e-10, 7.663061e-10, 
    1.329056e-09, -3.586251e-10, 5.04383e-09, 3.070056e-09, -6.501466e-10, 
    -5.802576e-10, -3.893661e-09, -1.975025e-10, -8.488996e-11, 
    -7.263701e-10, 8.581935e-11, -9.551826e-11, -3.155947e-10,
  1.064279e-09, 1.429612e-10, 4.542926e-10, -9.179644e-10, -2.696652e-09, 
    -1.840021e-10, -1.406437e-08, -1.855312e-09, 1.674721e-09, 1.78045e-09, 
    1.951719e-09, 5.862717e-09, -4.783942e-10, 1.447461e-09, 5.778759e-09, 
    5.056617e-10, -3.001497e-09, -3.110301e-09, -7.048797e-10, 7.797325e-09, 
    -4.906781e-09, -1.793751e-09, -8.85052e-10, 1.717808e-10, -1.866624e-09, 
    1.046476e-08, -1.949491e-08, -4.626543e-09, 3.759874e-08, -1.265477e-08, 
    -3.265751e-08, 1.082356e-09, -3.538048e-09, 7.853487e-10, 1.477304e-09, 
    -1.185367e-08, -1.393664e-09, -1.627498e-10, 3.800835e-09, 3.548417e-09, 
    1.613512e-09, -3.26088e-09, 8.472782e-09, -3.033215e-09, 1.13011e-08, 
    3.195964e-09, 1.863555e-09, 4.621626e-09, 7.224514e-09, -7.339231e-10, 
    1.601521e-09, 1.20923e-09, 6.204453e-09, -1.972239e-10, 7.678267e-09, 
    -6.187406e-11, 3.747402e-09, 6.501409e-10, -1.960598e-09, -1.474356e-08, 
    -4.061121e-09, 3.353762e-10, -1.961553e-09, -5.761342e-09, -6.406022e-10, 
    1.252067e-08, -8.915322e-10, 8.497182e-09, 1.061528e-08, -6.055245e-09, 
    -2.140894e-09, 3.416346e-09, -2.194213e-09, -1.604121e-10, 6.658143e-09, 
    4.928324e-11, -3.879421e-10, 1.844768e-09, 4.598192e-10, 1.272406e-08, 
    -3.690303e-09, -1.436879e-09, -5.232437e-11, -2.147544e-10, 5.359198e-10, 
    3.896901e-09, -7.670451e-10, -4.235972e-10, 1.412552e-09, 4.457377e-10, 
    1.260094e-08, 4.807919e-09, -5.976659e-10, -4.121117e-08, -1.531077e-09, 
    1.382244e-09, 4.943559e-10, -2.226159e-09, 8.536745e-10, -3.240984e-10, 
    8.611778e-11, 9.910472e-10, 8.762413e-11, 5.633751e-10, -2.789932e-09, 
    -3.568061e-10, 4.565095e-10, 1.140279e-09, -4.362164e-10, 5.358743e-09, 
    2.568811e-09, -3.713581e-10, -6.136816e-10, -4.068966e-09, 2.08729e-10, 
    -8.644747e-11, -8.64766e-10, 5.340439e-11, -9.312018e-11, -5.127276e-11,
  3.917535e-09, 4.081357e-10, -3.180958e-10, -9.345626e-10, -1.79358e-09, 
    -1.88686e-09, -2.350532e-09, -2.483887e-09, 4.271783e-10, 9.131895e-10, 
    -4.667982e-10, 4.984997e-09, -1.555179e-09, -1.238612e-08, 7.19325e-09, 
    5.442589e-10, -3.349379e-09, -5.705289e-09, -1.720835e-09, 1.000041e-08, 
    -1.598949e-09, -1.850083e-09, -8.740244e-10, 7.225367e-10, -1.520505e-09, 
    4.615117e-10, -1.199055e-08, -4.822027e-08, 1.936132e-08, -1.153995e-08, 
    -3.696334e-08, 1.054048e-09, -2.931415e-09, 5.401262e-10, 3.899856e-09, 
    -1.129195e-08, -2.141752e-09, -2.368097e-10, 9.059079e-09, 3.503692e-09, 
    6.728215e-10, -2.303807e-09, 1.351283e-08, -4.813426e-09, 7.677386e-09, 
    4.993694e-09, 2.022375e-09, 5.146219e-09, 1.264909e-08, -9.324665e-10, 
    3.24092e-09, 3.184482e-09, 7.933909e-09, -2.291586e-10, 9.038228e-09, 
    9.274004e-11, 6.284438e-09, 1.270712e-09, -3.581011e-09, -8.541555e-09, 
    1.652779e-09, 3.849266e-09, -1.962235e-09, -8.89337e-09, 5.920413e-09, 
    8.850122e-09, 4.814638e-11, 1.891846e-08, 1.055076e-08, -1.141075e-09, 
    -1.353612e-09, -7.22423e-10, -7.308927e-10, 3.549076e-09, 9.165774e-09, 
    -4.501999e-11, -5.410641e-10, 3.58439e-09, 4.768438e-10, 1.099176e-08, 
    -3.433286e-09, -5.313401e-09, -2.92772e-10, -2.108891e-10, 1.569106e-09, 
    4.009848e-09, -4.806566e-09, -7.180461e-10, 4.754622e-09, 5.476579e-10, 
    1.303619e-08, 1.068656e-09, -4.647376e-10, -2.301639e-08, 2.960405e-10, 
    2.217268e-09, -3.100126e-10, -1.267608e-08, 1.531873e-09, -8.015263e-10, 
    1.242029e-10, 9.197144e-09, -1.803286e-10, 8.161969e-10, -9.736993e-09, 
    -3.388038e-09, -9.679866e-10, -2.716149e-09, -3.916e-09, 9.614382e-09, 
    3.721425e-09, -8.649863e-10, 1.805006e-09, -4.873641e-09, -2.060176e-09, 
    -8.404299e-11, -7.265939e-10, 4.243716e-11, -8.756729e-11, 1.930403e-10,
  6.261928e-09, -2.500883e-09, -7.723884e-10, -2.768274e-10, -1.984972e-10, 
    -3.530715e-09, 3.342336e-09, -6.590597e-09, -1.770672e-10, 9.911219e-10, 
    -2.750937e-09, 2.942784e-09, 1.202238e-09, -1.022255e-08, 7.386802e-10, 
    -3.136904e-10, -4.125996e-09, -8.277027e-09, -2.813188e-09, 1.40231e-08, 
    2.193872e-09, -4.884612e-09, -8.192842e-10, 1.521528e-09, 1.157332e-10, 
    1.088551e-10, -2.990873e-08, -5.777758e-08, 1.044407e-08, -5.852996e-09, 
    -3.03998e-08, -7.661924e-10, -3.658783e-09, -1.571152e-10, 3.563741e-09, 
    -1.10698e-08, -2.757241e-09, -2.867253e-10, -9.263943e-09, 2.36551e-09, 
    -3.714445e-09, 4.181175e-09, 1.620938e-08, -8.310916e-09, 1.57408e-08, 
    1.970034e-08, 2.517709e-09, 2.770577e-09, 1.983269e-08, -1.200203e-09, 
    4.434774e-09, 1.801709e-09, 9.054526e-09, -4.571461e-10, 6.096639e-09, 
    2.341949e-10, 9.15378e-09, 1.958489e-09, -7.238413e-09, 3.914025e-10, 
    1.263226e-08, 6.079347e-09, -7.127596e-10, -6.163384e-09, 1.506646e-09, 
    6.067239e-09, 2.290165e-09, 4.281935e-08, 2.225954e-08, 9.053736e-09, 
    -4.780532e-11, 2.5178e-08, 6.547225e-10, 3.195112e-09, 1.194794e-08, 
    -1.792273e-10, -5.658691e-10, 7.608591e-09, 4.503391e-10, 1.700772e-08, 
    -1.850736e-09, -7.324637e-09, -1.736282e-10, -1.482817e-09, 3.267189e-09, 
    1.580474e-09, -6.396476e-09, -1.09344e-09, 8.673553e-09, 3.151911e-09, 
    6.160747e-09, -2.818865e-09, 1.061039e-09, 2.807091e-08, 1.007322e-09, 
    2.885076e-09, -4.900857e-09, -2.013439e-08, 2.86434e-09, -1.336377e-09, 
    1.1118e-09, 1.223139e-08, -5.830039e-10, 9.428014e-10, -2.597761e-08, 
    -2.061654e-09, 5.288882e-09, -9.947769e-09, 3.469893e-09, 1.390066e-08, 
    4.522633e-09, -3.597734e-09, 2.943239e-09, -5.880111e-09, -8.651625e-09, 
    -6.511982e-11, -5.359482e-10, 4.802025e-11, -3.903722e-11, 1.073147e-09,
  8.185509e-09, -5.170136e-09, -1.061494e-09, -9.614496e-10, 5.153993e-10, 
    -2.865136e-09, -5.441052e-10, -1.906369e-08, -1.892886e-10, 1.163301e-09, 
    -1.492367e-09, -7.808012e-10, 6.099867e-10, -5.500738e-10, -9.055725e-10, 
    1.124391e-09, -6.643762e-09, -8.37295e-09, -3.096368e-09, 1.806563e-08, 
    3.794185e-09, -9.920939e-09, -5.673542e-10, 1.480373e-09, 7.218546e-10, 
    1.105036e-10, -1.40293e-08, -5.05749e-08, 1.254114e-08, 7.288293e-09, 
    -3.067601e-08, -4.071524e-09, -5.084985e-09, -1.866056e-09, 1.278806e-09, 
    -1.312355e-08, -3.787113e-09, -2.721805e-10, -4.890035e-08, 4.927472e-10, 
    -1.214222e-08, 9.717894e-09, 1.591062e-08, -1.383427e-08, 2.475468e-08, 
    3.833503e-08, 5.225473e-09, -4.663576e-10, 2.978592e-08, -1.5323e-09, 
    4.542819e-09, -3.593755e-09, 8.367572e-09, -1.263811e-09, 4.468073e-09, 
    3.944649e-10, 9.640587e-09, 9.842666e-10, -1.163845e-08, 1.054882e-08, 
    5.612833e-09, 5.184631e-09, 4.163212e-10, -2.776119e-09, -2.612615e-09, 
    7.130041e-09, 1.221764e-08, 5.631051e-08, 2.349435e-08, 1.433153e-08, 
    -2.33581e-09, 3.055101e-08, -9.164864e-09, -2.442562e-10, 1.38161e-08, 
    -3.215064e-10, -6.61494e-10, 1.502528e-08, 3.198096e-10, 2.814744e-08, 
    -2.106447e-09, -4.414961e-09, 2.212346e-10, 1.120782e-09, 4.629442e-09, 
    -3.639116e-10, -5.329866e-09, -2.127308e-09, 4.13138e-09, 7.792835e-09, 
    6.623395e-10, -2.788772e-09, 2.605262e-09, 7.991484e-08, -9.167707e-10, 
    3.242258e-09, -1.302758e-08, -3.001787e-09, 5.04906e-09, -1.982062e-09, 
    1.152557e-09, 3.628429e-09, -7.283312e-10, 5.210552e-10, -9.709368e-09, 
    3.006221e-09, 1.936655e-10, -6.989069e-09, 1.23016e-08, 1.434853e-08, 
    2.745594e-09, -8.467566e-09, -1.62629e-10, -6.715652e-09, -1.121469e-08, 
    -2.925731e-11, -1.537046e-10, 6.150103e-11, 1.28253e-12, 2.259469e-09,
  5.396828e-09, -4.310948e-09, -2.619913e-10, -4.088747e-10, -1.317574e-09, 
    2.719958e-10, -5.14882e-09, -2.639575e-08, -1.13198e-09, -1.336218e-09, 
    4.460503e-10, -4.516323e-09, 3.845003e-09, 1.291221e-08, 6.83508e-09, 
    1.806512e-09, -1.120375e-08, -6.430014e-09, -3.072273e-09, 2.009517e-08, 
    8.681297e-09, 3.422429e-09, -5.635172e-09, 6.589289e-10, 1.610488e-09, 
    3.760761e-10, 5.669233e-08, -3.559273e-08, 5.588902e-09, 1.806171e-08, 
    -3.595346e-08, -5.187133e-09, -6.535458e-09, -3.511843e-09, 4.075673e-10, 
    -1.582254e-08, -5.623002e-09, -9.902834e-11, -8.155394e-08, 
    -1.176113e-09, -2.493702e-08, 1.147163e-08, 1.517861e-08, -2.263552e-08, 
    7.039665e-08, 4.011014e-08, 9.537473e-09, -2.86137e-09, 4.168288e-08, 
    -1.985686e-09, 1.823558e-09, -1.168968e-08, 8.047072e-09, -5.901142e-10, 
    7.070125e-09, 4.75211e-10, 4.67702e-09, -1.248964e-10, -1.329881e-08, 
    1.090068e-08, -1.010847e-08, 3.24809e-09, 2.012143e-09, -2.382433e-09, 
    -3.754337e-09, 1.026513e-08, 1.637051e-08, 4.302905e-08, 2.235544e-08, 
    1.318909e-08, -5.864422e-09, 4.120869e-08, -1.371433e-08, -1.918295e-09, 
    1.469633e-08, -5.127845e-10, -5.708287e-10, 2.446191e-08, -5.885852e-11, 
    2.910133e-08, -3.96318e-09, -6.929845e-09, 8.700169e-10, 4.54861e-10, 
    -2.051138e-09, -1.210992e-09, -9.041457e-09, -2.636114e-09, 
    -2.280117e-09, 6.545577e-09, -1.36896e-09, -1.230796e-09, 3.809944e-09, 
    9.704414e-08, -4.150024e-09, 3.398441e-09, -1.988301e-08, 8.854329e-09, 
    7.715016e-09, -2.608306e-09, 8.265602e-10, -1.030383e-09, -1.385292e-09, 
    -6.069776e-10, 1.054315e-08, 6.467644e-10, -7.894357e-09, 3.972104e-09, 
    1.44646e-08, 6.522384e-09, 1.05689e-09, -1.045413e-08, -6.522782e-10, 
    -7.129643e-09, -1.365572e-08, -1.844e-11, 5.767475e-11, 7.057643e-11, 
    5.361755e-11, 3.701302e-09,
  1.479634e-09, -5.070433e-10, -9.879386e-10, 3.677599e-09, -2.403794e-09, 
    2.588479e-09, -6.392952e-09, -1.618002e-08, -8.421239e-09, -6.115272e-09, 
    -2.605759e-09, -3.373714e-09, 6.45889e-09, 7.079507e-09, 9.525138e-09, 
    -8.023058e-10, -1.396475e-08, -2.67562e-09, -3.439098e-09, 2.002054e-08, 
    4.637798e-09, 3.028845e-09, -6.188543e-09, -1.902265e-09, 2.514071e-09, 
    5.868515e-10, 8.254972e-08, -1.904471e-08, -6.146314e-08, 2.320155e-08, 
    -3.192611e-08, -9.526048e-09, -8.823235e-09, -7.203312e-09, 
    -1.138574e-10, -1.576126e-08, -5.30049e-09, 2.07649e-10, -8.744348e-08, 
    5.247319e-09, -4.260669e-08, 4.640526e-09, 1.492995e-08, -3.167595e-08, 
    2.631691e-08, 3.151229e-08, 8.758491e-09, -4.106198e-09, 5.268813e-08, 
    -2.483727e-09, -7.811352e-10, -1.064376e-08, 1.161493e-09, -1.898593e-09, 
    8.694154e-09, 4.310436e-10, -8.381903e-09, 5.29509e-09, -1.105829e-08, 
    -5.804573e-09, 4.424749e-09, 2.549086e-09, 3.327614e-10, -1.637727e-09, 
    -3.348089e-09, 3.468324e-08, 2.708202e-08, 4.592323e-08, 2.143611e-08, 
    5.125798e-09, -4.440614e-08, 7.568366e-08, -9.609892e-09, -2.664706e-09, 
    1.628153e-08, -9.289352e-10, -1.160572e-09, 3.109203e-08, -1.168101e-09, 
    1.747907e-08, -2.742297e-09, -1.165328e-08, 1.651841e-09, 6.913297e-10, 
    -2.77214e-09, -1.578769e-09, -1.204262e-08, -6.208438e-10, -2.718942e-08, 
    3.226e-08, -2.386287e-10, -1.721423e-09, 4.713741e-09, 7.106792e-08, 
    -5.668255e-09, 3.08076e-09, -1.845617e-08, 2.071226e-08, 9.954078e-09, 
    -2.83369e-09, 3.323066e-10, -8.778294e-10, -1.37166e-09, -1.575323e-09, 
    -4.956348e-09, -5.274103e-09, -6.115215e-10, 8.9683e-09, 6.342987e-09, 
    7.156586e-10, -2.991101e-09, -5.251877e-09, -2.901288e-10, -6.208495e-09, 
    -2.025814e-08, -8.649863e-11, 5.153353e-10, 4.441425e-11, 8.395773e-11, 
    6.210314e-09,
  -6.62908e-10, -2.484057e-11, -3.586365e-09, 2.307792e-08, -1.086335e-09, 
    2.01203e-09, -5.204811e-09, 4.128026e-09, -2.453345e-08, -1.217626e-08, 
    -4.558444e-09, 2.831939e-09, 2.373099e-09, 3.233311e-09, 1.631429e-08, 
    -1.222153e-08, -1.738668e-08, 3.526111e-09, -3.111992e-09, 1.627603e-08, 
    1.050012e-09, 1.098613e-09, -1.27045e-10, -7.621793e-09, 3.327557e-09, 
    -9.310952e-11, 4.721096e-08, -8.921006e-09, -6.494651e-08, 1.888765e-08, 
    -2.400407e-08, -4.552533e-09, -1.954123e-08, 9.798896e-09, -2.92232e-10, 
    -1.101949e-08, -2.125995e-09, 8.625491e-10, -7.15346e-08, 2.201053e-08, 
    -6.331963e-08, 4.029459e-09, 1.356483e-08, -4.042559e-08, 3.065355e-08, 
    1.593452e-08, 2.382876e-10, -2.95978e-09, 4.848777e-08, -2.924594e-09, 
    -3.614957e-09, -5.654726e-09, -1.641128e-08, -1.081298e-09, 9.64074e-09, 
    1.873559e-10, -3.131385e-08, 1.060778e-08, -2.41958e-09, -1.561958e-08, 
    2.171413e-08, 4.665139e-09, 5.957759e-10, 1.128148e-09, -3.018011e-09, 
    1.789774e-07, 1.128403e-07, 6.158592e-08, 2.952879e-08, -2.483148e-08, 
    -6.056854e-08, 2.806991e-08, -4.423157e-09, -4.027186e-09, 2.061717e-08, 
    -1.201329e-09, -1.191928e-09, 3.530742e-08, -3.358837e-09, 2.931415e-09, 
    -5.423544e-09, -1.761599e-08, 2.419966e-09, 5.678658e-10, -3.369109e-09, 
    -7.640722e-09, -4.521382e-09, 3.034188e-09, -5.895009e-08, 4.502058e-08, 
    7.261747e-10, 7.647463e-09, 4.452531e-09, 3.368594e-08, -1.052121e-08, 
    1.934279e-09, -8.78756e-09, 4.993393e-08, 9.553787e-09, -3.176285e-09, 
    -4.000071e-10, 2.56227e-09, 2.573792e-09, -3.414563e-09, -1.840561e-08, 
    -8.326822e-09, 1.251919e-09, 5.173888e-09, 2.749971e-09, -1.498563e-09, 
    -7.146525e-09, 4.564527e-11, -9.237056e-10, -4.453511e-09, -1.222372e-08, 
    -2.770946e-10, 3.28896e-10, 2.007994e-10, 1.126033e-10, 8.046584e-09,
  -3.644232e-09, -8.615189e-10, 7.68523e-11, 4.630442e-08, 1.730143e-09, 
    3.655714e-09, -2.532317e-09, 9.684015e-09, -3.426067e-08, -1.182184e-08, 
    -9.51843e-10, 7.875371e-09, 6.491518e-11, 1.33582e-10, 1.203483e-08, 
    -9.548449e-09, -2.43445e-08, 1.060931e-08, 4.202789e-10, 7.29051e-09, 
    1.1363e-09, 5.940478e-09, 3.690843e-10, -1.423473e-09, 2.116508e-09, 
    -2.180514e-09, 1.373184e-08, -8.257814e-09, 5.887273e-10, 7.565006e-09, 
    -1.646072e-08, -4.184642e-09, -1.962076e-08, 4.19621e-08, 2.693525e-09, 
    9.721361e-10, 1.146083e-09, 2.060503e-09, -3.904421e-08, 5.441914e-08, 
    -7.653327e-08, 5.249376e-09, 1.188879e-08, -4.384544e-08, 2.356893e-08, 
    1.643218e-08, -9.633482e-09, -8.093565e-09, 3.918711e-08, -3.530225e-09, 
    -6.623068e-09, -2.229706e-08, -3.922095e-08, 1.204592e-09, 1.478838e-08, 
    1.948308e-10, -6.257534e-08, 1.06838e-08, 1.608509e-08, 1.144187e-09, 
    7.002882e-09, 3.250307e-09, 1.809497e-09, 8.294421e-09, -1.290865e-08, 
    1.707041e-07, 1.483635e-07, 2.68596e-08, 3.142844e-08, -3.345929e-08, 
    -4.955922e-08, 4.421759e-08, -1.567861e-08, -4.001208e-10, 2.935219e-08, 
    -8.807888e-10, 1.069381e-09, 4.24467e-08, -5.541898e-09, -6.724008e-10, 
    -6.96636e-09, -2.772926e-08, 4.062429e-09, -1.154262e-09, 3.765763e-09, 
    -8.670725e-09, -3.043795e-09, 5.258983e-09, -5.409166e-08, 3.654085e-08, 
    8.837446e-10, 2.192462e-08, 3.331209e-09, 6.842122e-09, -2.30466e-08, 
    3.155321e-10, 3.487571e-10, 8.352879e-08, 8.654354e-09, -5.084325e-09, 
    8.618599e-10, 1.626347e-09, 6.744056e-09, -5.584951e-09, -1.92407e-08, 
    -9.412702e-09, -5.607831e-09, -2.229001e-09, 4.258311e-09, -3.624564e-09, 
    -8.610471e-09, 2.54812e-09, -1.162789e-09, -3.049024e-09, 4.430376e-09, 
    -4.691685e-10, 6.970424e-12, 1.802061e-10, 1.444143e-10, 7.786639e-09,
  -5.199354e-09, 2.828642e-09, 2.389129e-09, 7.830829e-08, 7.425683e-09, 
    1.113551e-08, -1.376179e-09, 4.152071e-09, -1.98844e-08, -4.493813e-09, 
    2.902993e-09, 6.43513e-09, -2.058073e-09, -4.184471e-09, 1.027729e-09, 
    1.994196e-08, -3.859861e-08, 1.813544e-08, 6.670859e-09, 2.42153e-11, 
    1.974354e-08, -1.100591e-08, -2.873981e-08, 9.399628e-10, -3.346713e-09, 
    -6.87146e-09, -4.738467e-10, -1.120679e-08, -1.603132e-08, -6.537448e-09, 
    -1.541048e-08, 1.611647e-08, -1.192359e-08, 5.901416e-08, 2.25873e-09, 
    9.598125e-09, 4.381172e-09, 4.188095e-09, 8.998904e-08, 1.041009e-07, 
    -7.137237e-08, 5.240963e-09, 1.56509e-08, -4.175127e-08, -9.915198e-09, 
    -2.874413e-08, -1.61121e-08, 1.318409e-08, 2.839454e-08, -4.708468e-09, 
    -8.687422e-09, -5.916627e-08, -7.587799e-08, -1.602757e-10, 2.358428e-08, 
    -3.052492e-11, -7.947301e-08, 4.371792e-09, 3.994661e-08, 1.977254e-08, 
    -2.32933e-09, 5.853735e-10, 2.917886e-09, 1.319611e-08, -4.043361e-08, 
    1.164466e-07, 1.132528e-07, -3.021e-09, 1.785588e-08, -1.715523e-08, 
    -1.613887e-08, 2.081855e-07, -3.672494e-08, 1.917556e-09, 3.370707e-08, 
    5.377387e-10, 2.152504e-09, 4.398154e-08, -8.121305e-09, -5.221636e-10, 
    -8.277539e-09, -3.592618e-08, 6.287053e-09, -5.396942e-09, 1.840488e-08, 
    -3.156401e-09, -3.691184e-09, 4.873414e-09, -4.192356e-08, 7.970755e-09, 
    5.452421e-10, 2.749327e-08, 1.446494e-09, -5.838147e-08, -4.512617e-08, 
    -9.255473e-10, 5.543598e-10, -4.72437e-09, 8.383495e-09, -9.395876e-09, 
    -1.352873e-11, -1.505434e-09, 4.126122e-09, -7.148444e-09, -2.25391e-08, 
    -2.33581e-08, -1.631042e-08, -1.17243e-08, 7.300741e-09, -3.277478e-09, 
    -7.541189e-09, 7.349854e-10, -4.673666e-10, -6.644996e-10, 6.296204e-09, 
    -6.91648e-10, -1.625011e-10, 2.462812e-10, 1.543441e-10, 5.426273e-10,
  -2.108317e-08, 6.545235e-09, 1.237282e-08, 1.212755e-07, 2.45854e-08, 
    1.672271e-08, -2.251284e-09, 2.563013e-09, 9.373196e-09, 4.650417e-09, 
    8.032487e-09, 3.227967e-09, -1.200476e-09, -1.004418e-08, 5.258016e-11, 
    5.087037e-08, -4.59441e-08, 2.972376e-08, -2.717472e-08, 4.70942e-09, 
    4.352438e-08, -9.485859e-09, -2.113899e-08, -3.083318e-08, -1.663335e-08, 
    -5.898926e-09, -5.100368e-07, -1.306324e-08, -1.814777e-08, 
    -2.219605e-08, -3.298868e-08, -4.4513e-08, -6.456975e-08, 6.193892e-08, 
    -2.682958e-08, 4.58511e-08, 1.102632e-08, 5.572076e-09, 1.337075e-07, 
    1.628744e-07, -5.958692e-08, 3.454318e-09, 1.75871e-08, -4.147641e-08, 
    -2.988605e-08, -1.600069e-07, -1.678546e-08, 6.183555e-08, 1.81779e-08, 
    -6.114895e-09, -7.004175e-09, -9.585978e-08, -1.098961e-07, 
    -2.693775e-09, 3.371927e-08, -1.183707e-09, -8.023113e-08, -3.163347e-09, 
    4.753767e-08, 3.419497e-08, 1.773685e-09, -2.518163e-11, 3.568232e-09, 
    1.529542e-08, -7.073921e-08, 3.297288e-08, 6.113981e-08, 1.110897e-08, 
    2.498217e-08, 4.549491e-08, 2.567896e-08, 2.325657e-07, -4.441046e-08, 
    2.440686e-09, 2.646467e-08, 2.952504e-09, 2.683592e-09, 3.999702e-08, 
    -1.056213e-08, 2.593765e-10, -8.33893e-09, -3.537255e-08, 7.981782e-09, 
    -6.147104e-09, 1.69444e-08, 8.338873e-09, 2.390829e-08, 2.793797e-09, 
    -3.908357e-08, -2.013837e-08, 4.499157e-10, 2.456394e-08, -3.682032e-10, 
    -1.705987e-07, -5.461931e-08, -9.209656e-10, -7.625601e-09, 3.11872e-08, 
    8.093991e-09, -1.411425e-08, 8.793677e-11, -9.296599e-10, -5.792579e-09, 
    -6.627928e-09, -5.339217e-08, -4.408747e-08, -3.462213e-08, -2.03284e-08, 
    1.360019e-08, -2.168406e-09, -5.596178e-09, -3.634739e-09, -2.499405e-10, 
    1.45593e-09, 1.40534e-09, -1.013063e-09, 7.173639e-11, 8.075673e-11, 
    1.232934e-10, -6.49203e-09,
  -3.369757e-08, 4.122057e-09, 7.718086e-09, 1.081884e-07, 2.197999e-08, 
    1.164062e-08, 2.031811e-09, 6.616574e-11, 2.405068e-08, 4.420713e-09, 
    4.589424e-09, -1.143803e-09, -3.875584e-09, -5.010099e-08, 4.638991e-09, 
    7.73102e-08, -4.23611e-08, 4.195454e-08, -3.787136e-08, 2.026877e-08, 
    3.161392e-08, -7.569497e-09, 2.895035e-09, -2.197453e-09, -2.731213e-09, 
    1.643571e-09, -4.900166e-07, -1.999729e-08, -1.444596e-08, -2.53533e-08, 
    -5.873778e-08, -4.507115e-08, -4.350181e-08, 8.687005e-08, -7.599704e-08, 
    1.20288e-07, 1.721603e-08, 6.745836e-09, 6.065613e-08, 2.287423e-07, 
    -7.146959e-08, 2.231786e-09, 1.555313e-08, -4.462519e-08, -1.272326e-08, 
    -1.7837e-07, -4.671847e-09, 1.221455e-07, 6.904202e-09, -7.182152e-09, 
    -5.280327e-09, -8.111158e-08, -1.514151e-07, -2.979141e-09, 4.062917e-08, 
    -4.057654e-09, -7.910671e-08, 5.565175e-09, 2.21902e-08, 5.420266e-08, 
    3.767468e-09, 7.958079e-13, 1.16305e-08, 1.542933e-08, -9.053506e-08, 
    -2.519221e-08, 1.894102e-08, 2.128979e-08, 3.721186e-08, 7.965821e-08, 
    2.82397e-08, 1.775616e-07, -3.713149e-08, 1.132298e-08, 2.707056e-08, 
    -3.111722e-09, 1.136669e-09, 3.322299e-08, -1.215512e-08, 1.396404e-08, 
    -7.617416e-09, -1.86242e-08, 1.064831e-08, -4.120807e-09, -6.635901e-10, 
    1.507578e-08, -6.858613e-09, 1.844455e-09, -3.994431e-08, -7.391463e-08, 
    1.009539e-10, 1.510682e-08, -7.613608e-10, -2.624413e-07, -2.968773e-08, 
    -2.594732e-09, -9.820791e-09, 4.652259e-08, 3.04135e-09, -1.749024e-08, 
    -2.159868e-08, 6.125305e-09, -1.092119e-08, -3.360405e-09, -4.368462e-08, 
    -6.763855e-08, -5.355582e-08, -2.102206e-08, 2.404602e-08, 4.150706e-10, 
    1.134595e-10, -3.964715e-09, 9.874839e-10, 1.073545e-09, -7.493099e-10, 
    -1.184503e-09, 1.22678e-09, -1.367937e-10, 7.546674e-11, 6.511982e-10,
  4.978943e-08, 1.281535e-09, 2.529532e-11, 4.90358e-08, 9.534517e-09, 
    8.224845e-09, 1.65266e-08, -7.219398e-09, 2.12803e-08, 4.702713e-09, 
    -2.810907e-10, -5.669506e-09, -3.381331e-09, -1.17769e-07, 6.305584e-09, 
    1.058888e-07, -3.987979e-08, 4.778633e-08, 8.38768e-08, 2.729013e-08, 
    -4.063679e-09, -6.044161e-10, 7.45132e-09, 2.157947e-09, 1.124334e-08, 
    5.081745e-09, -6.463137e-08, -2.180508e-08, -2.085727e-08, -2.950873e-08, 
    -7.222758e-08, -3.766701e-08, 6.528427e-08, 9.087859e-08, -1.108036e-07, 
    1.807394e-07, 2.217305e-08, 7.505946e-09, -2.742928e-08, 2.867498e-07, 
    -7.007253e-08, 5.341064e-09, 1.237157e-08, -5.028526e-08, -1.226653e-08, 
    -1.090208e-07, 2.612023e-08, 1.900355e-07, -8.269524e-09, -8.147545e-09, 
    -6.907172e-09, -5.222711e-08, -1.773093e-07, -4.285369e-09, 4.116406e-08, 
    -3.290552e-09, -7.38583e-08, -1.229011e-08, -1.279444e-08, 8.799788e-08, 
    3.118998e-10, -3.234391e-11, 5.404405e-08, 8.479458e-09, -9.690528e-08, 
    -5.110945e-08, -2.229791e-08, 2.254041e-08, 4.741725e-08, 1.488917e-08, 
    1.504026e-08, 2.254106e-07, -1.273776e-08, 1.322388e-08, 4.105598e-08, 
    -2.340511e-08, -1.515659e-09, 2.354409e-08, -1.239499e-08, 9.39288e-08, 
    -7.51271e-09, 8.478708e-09, 2.208299e-08, -4.029232e-09, -9.480743e-09, 
    4.401182e-07, -3.233636e-07, 1.014195e-08, -6.171129e-08, -1.308793e-07, 
    -1.123851e-09, -2.41448e-08, -6.925234e-10, -3.495564e-07, 2.691064e-08, 
    -5.270988e-09, -1.511556e-08, 1.761185e-08, 1.474461e-09, -2.080311e-08, 
    -4.67208e-08, 9.215178e-09, -1.72683e-08, -1.598153e-10, -9.080111e-09, 
    -1.067046e-07, -4.396003e-08, -2.327903e-08, 3.616645e-08, 6.099469e-09, 
    5.312188e-09, -2.043237e-09, 9.792416e-10, -7.15778e-09, -2.60826e-09, 
    -1.435421e-09, 3.287212e-09, -1.897398e-10, 1.250555e-11, 2.171811e-08,
  1.234952e-07, 6.134542e-10, -4.493131e-09, 6.442406e-09, -1.316835e-09, 
    8.671009e-09, 3.039372e-08, -7.605649e-09, 1.832746e-09, 7.457857e-11, 
    1.642775e-10, -3.422883e-09, -4.157641e-09, -8.847496e-08, 8.878715e-09, 
    1.028008e-07, -4.716559e-08, 5.444696e-08, 1.021129e-07, 2.592492e-08, 
    -2.441971e-08, -2.806019e-09, 2.985416e-09, -2.008505e-09, 8.662028e-09, 
    2.671641e-11, -4.25573e-08, -1.173532e-08, -4.418609e-08, -2.256604e-08, 
    -4.870321e-08, -2.789011e-08, 4.73616e-08, 4.0131e-08, -1.20247e-07, 
    1.99879e-07, 2.707285e-08, 8.287159e-09, -1.003123e-07, 3.391045e-07, 
    -1.303072e-08, 8.219672e-09, 1.44758e-08, -5.145509e-08, -4.217782e-09, 
    -8.115057e-08, 7.376661e-08, 2.677997e-07, -3.648684e-08, -1.047478e-08, 
    -4.282469e-09, -4.814058e-08, -2.022899e-07, -3.634068e-09, 3.766732e-08, 
    -2.295224e-09, -6.692835e-08, -1.59192e-08, -2.513538e-08, 1.259267e-07, 
    -3.076593e-09, -4.569074e-10, 1.026447e-07, -1.381943e-08, -8.325933e-08, 
    -3.07374e-08, -4.408469e-08, 2.070703e-08, 4.641629e-08, 7.164772e-09, 
    -2.785885e-08, 7.324581e-08, -1.687681e-09, 8.521965e-09, 4.96874e-08, 
    -8.49775e-09, -4.083319e-09, 1.148101e-08, -1.154082e-08, 1.549276e-07, 
    -3.15606e-09, 3.119776e-08, 3.879887e-08, 1.343437e-09, -7.837343e-09, 
    2.10128e-07, -2.203755e-07, 2.818695e-08, -6.029934e-08, -1.71087e-07, 
    -1.270337e-09, -1.531935e-07, -1.169894e-09, -4.346975e-07, 9.360747e-09, 
    1.005471e-08, 1.211936e-08, 1.023398e-08, 8.077677e-09, -2.50584e-08, 
    -6.163316e-08, -3.825619e-09, -1.01493e-08, 1.351587e-09, -2.128445e-09, 
    -7.738117e-08, -2.525951e-08, -2.502463e-08, 4.387061e-08, 1.937792e-08, 
    1.922558e-09, -6.131245e-09, -4.090225e-09, -1.86036e-08, -5.321454e-09, 
    -1.56482e-09, 4.09598e-09, -4.480007e-10, -6.472334e-11, 1.644787e-08,
  1.01266e-07, -1.014371e-09, -2.03151e-08, 1.790966e-09, 8.55988e-09, 
    2.315193e-08, 3.215945e-08, 3.249681e-09, -1.503912e-08, -4.74148e-09, 
    -3.475236e-09, -1.029434e-10, 5.634888e-10, 1.006034e-07, -1.333484e-08, 
    9.741364e-08, -4.612512e-08, 2.057999e-08, 1.582835e-08, -7.196945e-10, 
    -9.241774e-09, -1.194149e-08, 1.818705e-09, -2.023e-09, -6.028245e-10, 
    -4.264126e-08, -6.175981e-09, -5.455547e-09, -7.166312e-08, 1.153069e-09, 
    -1.364009e-08, -1.720497e-08, 1.06798e-08, 2.374424e-08, -9.476986e-08, 
    1.9285e-07, 3.05874e-08, 9.468295e-09, -1.136092e-07, 3.720957e-07, 
    8.110013e-08, 8.164022e-09, 2.351533e-08, -5.47478e-08, -2.322793e-09, 
    -1.043118e-07, 1.281692e-07, 3.172835e-07, -6.970683e-08, -1.241512e-08, 
    6.960192e-10, -4.83638e-08, -2.206018e-07, -2.483569e-09, 2.785457e-08, 
    -1.622425e-09, -7.570287e-08, -3.186293e-08, -1.723428e-08, 1.510234e-07, 
    -2.133731e-09, 1.753227e-08, 6.714998e-08, -4.582488e-08, -5.383714e-08, 
    -1.746201e-08, -5.236922e-08, 2.318637e-08, 3.702854e-08, 6.475886e-09, 
    5.256395e-07, -4.930308e-08, -2.321229e-08, 1.80209e-08, 4.811232e-08, 
    -9.43993e-09, -5.640999e-09, 1.024716e-09, -1.05735e-08, -2.307689e-08, 
    1.073943e-09, 5.471946e-08, 5.220232e-08, -6.79222e-10, -1.516185e-09, 
    4.369605e-08, 6.706642e-08, 3.785357e-08, -6.474068e-09, -1.902289e-07, 
    -5.84356e-09, -2.396399e-07, -2.571795e-09, -4.92802e-07, -1.099119e-08, 
    3.043716e-08, 2.914672e-08, 3.20054e-08, 2.305268e-08, -2.713685e-08, 
    -2.013286e-08, -2.702247e-08, -1.190325e-08, 1.121478e-09, -2.387759e-08, 
    -5.128737e-08, -4.578686e-08, -1.802579e-08, 4.281691e-08, 3.226324e-08, 
    -1.551825e-11, -9.947087e-09, -1.367556e-08, -2.540691e-08, 
    -3.859952e-09, -1.546914e-09, 3.270273e-09, -7.471606e-10, -1.003073e-10, 
    -8.844228e-08,
  7.712453e-08, -1.989804e-09, -1.069833e-08, -2.481727e-09, 1.494601e-08, 
    3.179565e-08, 3.975327e-08, 2.367807e-08, -2.27173e-08, 3.593925e-09, 
    -3.962555e-10, -1.969113e-09, -9.66719e-09, 1.088304e-07, 2.451145e-09, 
    8.260485e-08, -3.157048e-08, -1.178859e-08, -6.977314e-08, -4.914187e-08, 
    1.073732e-08, -2.101336e-08, 4.601191e-09, -7.102585e-10, -9.644793e-09, 
    -1.507427e-07, -1.614006e-08, -1.049654e-08, -9.483034e-08, 2.537894e-08, 
    4.99125e-09, -2.311668e-08, -2.098994e-08, 2.33959e-08, -6.415388e-08, 
    1.576532e-07, 2.944547e-08, 9.215739e-09, -1.252415e-07, 3.823488e-07, 
    1.511425e-07, 9.024404e-09, 2.646559e-08, -7.12125e-08, 4.764217e-09, 
    -1.204529e-07, 1.576549e-07, 3.221981e-07, -8.431228e-08, -1.303405e-08, 
    4.415881e-09, -5.741725e-08, -2.402729e-07, -7.107394e-09, 1.635625e-08, 
    -1.3722e-09, -9.859326e-08, -4.8482e-08, 3.141202e-09, 1.445976e-07, 
    3.245191e-10, 3.910105e-08, 2.683765e-08, -7.756881e-08, -3.997021e-08, 
    -1.575057e-08, -4.533928e-08, 1.415293e-08, 2.740563e-08, 2.970808e-09, 
    2.352218e-07, -7.791704e-08, -7.492741e-08, 3.279126e-09, 4.442001e-08, 
    -1.358029e-08, -7.784436e-09, -5.755084e-09, -9.946578e-09, -4.42372e-08, 
    2.623608e-09, 7.753069e-08, 5.252667e-08, -7.174089e-08, 1.927845e-09, 
    -2.140138e-08, 3.906865e-08, 3.540134e-08, 4.729259e-08, -1.663872e-07, 
    -1.242557e-08, -2.078011e-07, -4.983264e-09, -5.330041e-07, 
    -2.404198e-08, 3.757461e-08, 3.670754e-08, 3.237056e-08, 3.127485e-08, 
    -2.605296e-08, 4.179122e-08, -3.184406e-08, -1.687491e-08, 6.762662e-10, 
    -3.65149e-08, -1.022476e-07, -8.035323e-08, -1.182326e-08, 4.563384e-08, 
    3.207305e-08, -6.307914e-10, -1.327993e-08, -2.105463e-08, -2.5269e-08, 
    -1.600426e-09, -1.741148e-09, 2.472873e-09, -1.154262e-09, -1.140563e-10, 
    -7.074374e-08,
  6.562357e-08, -5.609877e-09, -2.420734e-09, -7.884978e-09, 6.993218e-09, 
    3.690855e-08, 5.454115e-08, 4.130186e-08, -1.404067e-08, -2.968932e-09, 
    9.416681e-10, -2.264403e-08, -4.48664e-08, -3.664616e-08, 2.581794e-08, 
    6.436598e-08, -2.061888e-08, 3.257594e-08, -6.159223e-08, -1.10498e-07, 
    1.310343e-08, 4.084961e-08, 1.091814e-08, 1.337526e-09, -3.402727e-08, 
    -2.140229e-07, -1.040542e-08, -5.470042e-09, -1.090206e-07, 1.969136e-08, 
    7.609401e-09, -3.7208e-08, -3.104435e-08, 1.525825e-08, -5.343315e-08, 
    1.24019e-07, 2.340678e-08, 8.350725e-09, -1.289164e-07, 3.676623e-07, 
    2.13298e-07, 1.169053e-08, 1.7763e-08, -8.442618e-08, 6.892492e-09, 
    -1.05748e-07, 1.433683e-07, 2.760017e-07, -7.473484e-08, -1.300788e-08, 
    6.851195e-09, -6.487574e-08, -2.680998e-07, -6.745381e-09, 5.741214e-09, 
    -8.112693e-10, -1.017739e-07, -9.896787e-08, 1.6986e-08, 1.257452e-07, 
    1.673584e-09, 4.056858e-08, -1.268921e-07, -8.779877e-08, -4.197588e-08, 
    7.161702e-09, -5.428547e-10, -5.161269e-09, 1.764113e-08, -8.238771e-09, 
    -2.852231e-07, -1.07536e-07, -6.779453e-08, -3.934815e-09, 4.747999e-08, 
    9.66736e-09, -1.46706e-08, -5.956451e-09, -9.120759e-09, -1.87971e-08, 
    1.909939e-09, 9.857812e-08, 4.973583e-08, -2.527626e-07, 2.887157e-08, 
    6.00711e-08, -5.167101e-08, 4.406877e-08, 1.02586e-07, -8.094128e-08, 
    -1.977014e-10, -1.440654e-07, -6.305356e-09, -5.478453e-07, 
    -6.814275e-09, 3.752718e-08, -1.445198e-08, 3.47269e-08, 4.461151e-08, 
    -2.240097e-08, 1.750392e-07, -1.537849e-08, -2.661693e-08, -1.045507e-09, 
    3.200887e-08, -1.05273e-07, -3.130651e-08, 3.670834e-09, 5.354343e-08, 
    2.59223e-08, -1.858439e-09, -1.211072e-08, -1.777028e-08, -2.094987e-08, 
    1.838316e-10, -2.036336e-09, 1.993357e-09, -1.143022e-09, -2.119833e-10, 
    -8.772361e-08,
  6.089061e-08, -1.607174e-08, 2.691365e-09, -1.351992e-08, -3.746948e-09, 
    3.848612e-08, 6.698195e-08, 6.744443e-08, 7.826145e-09, -4.16378e-10, 
    -9.603184e-09, -1.229601e-07, -3.642396e-08, -1.471765e-07, 4.896395e-08, 
    4.672966e-08, -3.541387e-08, 5.101543e-08, -6.030078e-08, 1.119283e-07, 
    1.829125e-08, 2.745616e-07, 7.784308e-09, 4.70834e-10, -1.823406e-08, 
    -8.704507e-08, -1.684913e-08, -5.779896e-09, -1.129411e-07, -7.00544e-09, 
    -7.988604e-09, -4.436885e-08, -2.587586e-08, 7.199168e-08, -4.924442e-08, 
    9.966942e-08, 1.414941e-08, 7.094627e-09, -1.174965e-07, 3.319842e-07, 
    3.944941e-07, -7.651693e-10, -7.307546e-08, -7.372969e-08, 7.362303e-09, 
    -5.587418e-08, 2.702848e-09, 2.036329e-07, -5.054204e-08, -1.153109e-08, 
    8.178802e-09, -9.730257e-08, -2.967425e-07, -2.08521e-09, 9.341192e-10, 
    -1.265903e-10, -6.367833e-08, -1.512061e-07, 1.385537e-08, 1.445399e-07, 
    1.399656e-09, -1.479049e-08, -1.322836e-07, -8.176603e-08, -5.005315e-08, 
    -1.804722e-09, 2.05452e-08, -2.288749e-08, 1.959933e-08, -3.049792e-08, 
    -3.617325e-07, -2.529629e-08, -2.569988e-08, 5.211803e-09, 3.335743e-08, 
    2.416476e-08, -7.956942e-09, -2.855813e-09, -7.57027e-09, -7.196746e-08, 
    -2.848424e-10, 1.019108e-07, 4.244538e-08, -1.072397e-07, 6.321164e-08, 
    -6.170978e-09, 1.496332e-07, 8.232581e-08, 1.39761e-07, 5.811427e-08, 
    -8.444715e-09, -1.123252e-07, -5.984305e-09, -5.294775e-07, 5.939972e-08, 
    1.439021e-07, -1.489065e-07, 7.695479e-08, 6.253134e-08, -1.512636e-08, 
    2.244712e-07, -3.012332e-09, -3.092936e-08, -3.915019e-09, 4.045859e-08, 
    -3.919632e-08, 2.923497e-08, 2.270571e-08, 4.826751e-08, 1.480447e-08, 
    3.73069e-09, -3.975913e-09, 1.233445e-09, -2.054304e-08, -1.85139e-10, 
    -2.775766e-09, 5.953325e-09, -1.238398e-09, -5.414194e-10, -1.509671e-07,
  5.327615e-08, -3.397076e-08, 1.141416e-10, -1.107105e-08, -1.282501e-08, 
    3.920331e-08, 6.405958e-08, 6.590199e-08, 1.975855e-08, -2.016805e-09, 
    4.210733e-09, -1.812891e-07, 1.102558e-08, -9.846462e-08, 1.936064e-08, 
    2.802317e-08, -4.795599e-08, 3.439209e-08, -4.917513e-08, -8.535244e-08, 
    2.415375e-07, 1.532085e-07, -3.143368e-07, -1.046849e-07, -1.628769e-08, 
    -2.9082e-08, -2.863294e-08, -7.583594e-09, -1.176497e-07, -3.064065e-08, 
    -1.523949e-08, -5.142442e-08, -1.837634e-08, 4.653953e-08, -4.149138e-08, 
    7.686344e-08, -9.957375e-10, 5.538993e-09, -1.033807e-07, 2.858911e-07, 
    2.875734e-07, -3.637656e-07, -9.574558e-08, -7.572038e-08, 6.523805e-09, 
    -1.278295e-09, -6.188179e-08, 1.325774e-07, -4.094831e-08, -9.506422e-09, 
    8.602427e-09, -1.714593e-07, -3.193269e-07, 1.355993e-08, -6.498402e-09, 
    -1.682565e-10, -4.701792e-08, -1.509744e-07, -5.421953e-09, 1.831979e-07, 
    -8.051302e-10, -9.787482e-08, -6.538562e-08, -5.349999e-08, 
    -7.535181e-08, -3.017658e-08, 1.672561e-08, -3.203058e-08, 2.283446e-08, 
    -4.27633e-08, -2.83901e-08, -1.285557e-07, -9.701125e-09, 1.646185e-09, 
    3.112491e-08, 4.048138e-08, 3.327358e-09, -1.677677e-09, -8.110424e-09, 
    -5.538527e-08, 2.171646e-09, 9.329538e-08, 3.147079e-08, -3.599826e-08, 
    8.417032e-08, -1.617855e-08, 4.161304e-07, 9.390783e-08, 1.788023e-07, 
    1.710858e-07, -4.996946e-08, -1.083357e-07, -4.52178e-09, -5.025879e-07, 
    1.243855e-07, 6.34637e-08, -1.916424e-07, 3.057012e-07, 7.712879e-08, 
    -3.355872e-08, -4.453045e-08, 5.591247e-09, -2.576394e-08, -5.990898e-09, 
    6.491064e-09, -9.714086e-09, 4.278536e-08, 3.935202e-08, 3.128298e-08, 
    -1.421995e-09, 2.067873e-08, -1.130957e-09, 1.732747e-08, -2.636921e-08, 
    -1.845819e-09, -3.473838e-09, 1.040362e-08, -1.344944e-09, -8.165131e-10, 
    -5.717766e-08,
  4.363204e-08, -5.571241e-08, -3.846594e-10, -1.456272e-09, 3.811294e-09, 
    2.557709e-08, 4.188638e-08, 4.136695e-08, 2.457165e-08, 1.383142e-08, 
    3.197187e-08, -2.955477e-08, 4.334146e-08, -4.185205e-08, -1.273705e-07, 
    4.197341e-08, -7.160423e-08, 2.357848e-08, -2.77178e-08, -7.868101e-08, 
    8.414889e-08, 1.879056e-08, -8.729143e-08, 4.198142e-08, -1.846445e-09, 
    -4.442569e-08, -4.897987e-08, -6.61845e-09, -1.166797e-07, -5.480234e-08, 
    1.043678e-07, -1.074119e-08, -2.748897e-08, 5.183068e-08, 2.784731e-08, 
    5.534633e-08, -2.115686e-08, 5.522139e-09, -9.181127e-08, 2.357616e-07, 
    2.157535e-07, 6.170734e-08, -9.491114e-08, -8.29104e-08, 1.52346e-09, 
    1.840664e-08, -8.105189e-09, 7.401235e-08, -2.784608e-08, -4.575767e-09, 
    8.769291e-09, -3.032569e-07, -3.271157e-07, 1.172347e-08, -1.358935e-08, 
    -7.607525e-09, -2.756514e-08, -1.185897e-07, -2.724919e-08, 1.828793e-07, 
    -4.048559e-09, -1.366311e-07, 1.403083e-08, -2.51529e-08, -1.283818e-07, 
    -4.111001e-08, -2.780718e-08, -3.366875e-08, 1.564314e-08, -4.108909e-08, 
    -5.654164e-08, -1.899508e-07, -1.287134e-08, -3.510735e-08, 3.521551e-08, 
    2.352823e-08, -7.873808e-09, 1.475996e-09, -3.219662e-09, -8.337162e-08, 
    -3.424532e-09, 8.915241e-08, 1.556788e-08, -4.133818e-08, 7.428554e-08, 
    -3.882377e-08, 4.940211e-07, 4.123393e-08, 2.031098e-07, 2.571338e-07, 
    -1.18296e-07, -1.129842e-07, -9.713887e-09, -4.395226e-07, 1.570446e-07, 
    -1.931486e-07, -2.659853e-07, 2.827124e-08, 8.610397e-08, -5.492383e-08, 
    2.291989e-08, 6.802239e-10, -1.764647e-08, -5.117016e-09, 4.249029e-08, 
    -4.573104e-08, -2.929727e-08, 1.024802e-08, 1.183258e-08, -1.670043e-08, 
    -2.357064e-08, -4.881196e-08, 4.899505e-09, -2.071312e-08, 1.200982e-08, 
    -3.531102e-09, 1.044063e-08, -1.450278e-09, -8.897487e-10, 1.19968e-09,
  4.102401e-08, -8.846666e-08, 7.336098e-09, 1.326464e-08, 2.438958e-08, 
    1.073897e-08, -9.060955e-09, -1.361866e-08, 1.15075e-08, 4.211608e-08, 
    3.064883e-09, 2.85678e-08, 5.033939e-09, -8.00685e-09, -2.64473e-07, 
    6.279352e-08, -8.856466e-08, 2.138472e-08, -2.999653e-08, -2.727916e-09, 
    -7.634947e-08, -5.550157e-08, -2.991248e-08, -2.877857e-08, 6.113044e-08, 
    -6.330936e-08, -2.295826e-08, -6.480491e-09, -1.142613e-07, 
    -7.565393e-08, 2.072226e-07, 1.432113e-09, -2.353784e-08, 6.659332e-08, 
    2.508898e-08, 2.402237e-08, -4.781932e-08, 7.562392e-09, -6.896551e-08, 
    1.508814e-07, 8.104551e-08, 2.213504e-07, -2.784986e-08, -8.398007e-08, 
    -2.048068e-09, 9.151677e-09, 1.949812e-07, 4.05023e-08, -2.297527e-08, 
    2.717115e-11, 9.228074e-09, 1.140778e-07, -3.044993e-07, 8.226266e-09, 
    -1.865048e-08, -1.082071e-08, -2.303193e-08, -8.615697e-08, 4.51629e-08, 
    1.334643e-07, -4.45732e-09, -7.642041e-08, 3.222578e-08, 7.219043e-09, 
    -1.941175e-07, -4.07e-08, -2.245122e-08, -2.454669e-08, 4.882054e-09, 
    -2.207537e-08, -7.158872e-08, -2.04814e-07, -3.513412e-08, -7.968436e-08, 
    2.211409e-08, 6.847927e-09, -3.481071e-08, 2.195861e-10, -1.031461e-08, 
    -9.317785e-08, -7.662265e-09, 9.880697e-08, -1.79341e-09, -9.314874e-08, 
    4.159835e-08, -1.096134e-08, 3.65951e-07, -1.065143e-08, 2.004833e-07, 
    3.249504e-07, -8.815721e-08, -1.196844e-07, 5.855327e-09, -3.185273e-07, 
    -6.239281e-08, -2.918493e-07, -1.782687e-07, -6.804714e-08, 9.235771e-08, 
    -6.477352e-09, 1.238561e-08, 2.102873e-08, -1.08945e-08, 2.996003e-09, 
    1.380954e-09, -5.73192e-08, -9.160055e-08, -1.394062e-08, -8.750135e-09, 
    -2.69257e-08, -1.629076e-08, -4.893911e-08, -5.172649e-08, 6.720597e-09, 
    7.160145e-08, -2.927709e-09, 9.631918e-09, -3.055803e-09, -8.74266e-10, 
    -2.677041e-08,
  1.2171e-07, -1.316486e-07, 1.67434e-08, 3.186443e-08, 4.476425e-08, 
    1.638529e-08, -1.818364e-07, -1.243204e-07, -6.59719e-09, -5.99411e-08, 
    1.16113e-07, 2.238301e-07, -7.063221e-08, -1.153391e-07, -2.638685e-07, 
    6.388512e-08, -1.026312e-07, 2.308201e-08, -3.0064e-08, 3.501287e-08, 
    -6.949307e-08, -6.400222e-08, -1.775214e-08, -6.148429e-08, 2.379373e-07, 
    -5.466103e-08, -2.218889e-08, -9.403664e-09, -1.136295e-07, 
    -7.991952e-08, 7.963496e-08, -6.931884e-09, -1.70009e-08, 5.442308e-08, 
    2.231656e-08, -4.263882e-09, -7.610278e-08, 1.060113e-08, -4.58885e-08, 
    6.883782e-08, 1.111232e-09, 7.834439e-08, 4.456638e-09, -8.046771e-08, 
    -2.225704e-09, -6.90369e-09, 2.976441e-07, 1.888213e-08, -2.125997e-08, 
    3.257739e-09, 8.991918e-09, 1.947192e-07, -2.360479e-07, 1.49064e-08, 
    -2.389049e-08, -2.641514e-10, -3.84245e-08, -7.267671e-08, 3.968481e-08, 
    1.533007e-08, 1.691484e-08, 3.996166e-08, 1.198858e-07, 2.420794e-08, 
    -2.367984e-07, -3.401846e-08, 8.428799e-09, -2.15793e-08, -2.531976e-09, 
    4.577089e-09, -8.094611e-08, -1.970947e-07, -8.041997e-08, -8.25591e-08, 
    1.643622e-08, 2.09053e-09, -2.592236e-08, 6.039045e-10, -2.025696e-08, 
    -1.940227e-07, -8.116956e-09, 1.128824e-07, -3.323777e-08, -7.87133e-08, 
    9.398451e-08, -2.621795e-08, 1.84595e-07, -1.691654e-08, 2.062147e-07, 
    3.367995e-07, 5.47596e-08, -1.209962e-07, 8.1655e-09, -1.885817e-07, 
    -1.6334e-07, -3.213519e-07, -4.063953e-08, -4.101406e-08, 6.732699e-08, 
    -2.379636e-09, 2.751955e-08, 1.145157e-07, -5.823637e-09, 7.030621e-09, 
    3.488464e-08, -2.914379e-08, -1.688122e-07, -2.445967e-08, -2.669043e-08, 
    -3.360418e-08, -2.513542e-08, 1.104428e-08, -3.490749e-08, 7.107758e-09, 
    4.472651e-08, -1.951923e-09, 9.263715e-09, -3.42304e-09, -8.677432e-10, 
    -2.876635e-08,
  1.235127e-06, -1.502616e-07, 2.359752e-08, 3.127138e-08, 3.716161e-08, 
    5.744153e-08, -3.806185e-07, -2.660242e-07, -9.902806e-08, -2.697175e-08, 
    1.907756e-08, 1.675538e-07, -7.294113e-08, -2.861598e-07, -1.388071e-07, 
    6.22782e-08, -1.354027e-07, 4.89182e-08, -3.013376e-08, -3.007665e-08, 
    -3.198761e-08, -5.369623e-08, -3.630464e-08, -3.513082e-08, 
    -2.513048e-09, -2.925617e-08, -4.356389e-08, -8.583243e-09, 
    -1.066029e-07, -8.891936e-08, -7.477183e-08, -1.170952e-08, 
    -2.748845e-08, 3.868843e-08, 7.533038e-08, 2.003162e-09, -9.780418e-08, 
    1.247378e-08, -3.477987e-08, -8.368147e-09, 7.562971e-08, 7.467361e-08, 
    -1.629692e-08, -6.946988e-08, 4.093863e-10, 4.900812e-09, 2.171288e-07, 
    5.95702e-09, -2.072936e-08, 3.967578e-09, 8.315823e-09, -9.327414e-08, 
    -2.021715e-07, 2.194117e-08, -3.138122e-08, -1.043759e-09, 5.474362e-09, 
    -9.879597e-08, 1.100935e-08, 2.643361e-08, 1.713556e-08, -4.260676e-08, 
    2.704444e-07, 6.160931e-08, -2.483816e-07, -2.768786e-08, 3.350613e-08, 
    -2.171805e-08, -1.058913e-08, 7.769245e-09, -7.713561e-08, -1.735121e-07, 
    -7.146286e-08, -9.238738e-08, 1.208916e-08, -1.086732e-09, -1.240522e-08, 
    2.132026e-09, -1.755143e-08, -1.261197e-07, -5.201628e-09, 1.307389e-07, 
    2.204882e-08, -6.090261e-08, 9.74062e-08, -2.889044e-08, 2.81799e-08, 
    -1.041906e-08, 2.091692e-07, 3.185466e-07, -4.908543e-08, -1.288432e-07, 
    1.053024e-10, -5.580051e-08, -2.076011e-07, -2.796477e-07, -4.984049e-08, 
    -1.735316e-08, 6.751031e-08, 1.622079e-08, 9.235009e-09, 5.070474e-08, 
    -3.833968e-09, 7.16414e-09, -3.021194e-08, 9.418727e-09, -2.002253e-07, 
    -2.990191e-08, -3.908963e-08, -5.032757e-08, -2.81143e-08, 7.623839e-10, 
    1.00938e-08, 3.052492e-09, 7.200015e-09, -5.993684e-10, 7.497576e-09, 
    -3.10542e-09, -7.468799e-10, -2.513775e-08,
  1.035514e-06, -9.696242e-08, 3.53063e-08, 1.907352e-08, 8.468379e-08, 
    -4.952602e-08, -1.061192e-07, -5.189935e-08, -5.546741e-08, 3.4957e-09, 
    -3.854467e-08, 1.092605e-07, -6.547867e-08, -3.150791e-08, -2.653206e-08, 
    6.696579e-08, -1.828992e-07, 1.766807e-08, -7.699654e-09, -1.178504e-07, 
    4.089372e-09, -4.45562e-08, 6.31548e-08, -2.266046e-08, -1.39493e-07, 
    -1.841028e-08, -5.260739e-08, -6.437688e-09, -1.020003e-07, -9.40118e-08, 
    -9.150818e-08, 2.152041e-08, -5.083933e-08, 1.832012e-08, 1.106156e-07, 
    8.395148e-09, -1.111202e-07, 1.262171e-08, -2.559824e-08, -5.96425e-08, 
    1.072507e-07, 2.823801e-07, -5.103004e-09, -5.780175e-08, -1.355431e-09, 
    -7.145843e-09, 1.083142e-07, 1.186149e-08, -3.005192e-08, 3.336666e-09, 
    7.312863e-09, -1.575965e-07, -1.744068e-07, 2.643889e-08, -3.997248e-08, 
    -1.554326e-09, 2.479902e-08, -1.857076e-07, -2.40702e-09, 9.665534e-08, 
    1.448324e-07, -3.385668e-08, 5.053396e-07, 1.354351e-07, -2.252614e-07, 
    -2.578264e-08, 2.711414e-08, -2.777887e-08, -2.146118e-08, -7.852918e-10, 
    -8.029286e-08, -1.512834e-07, -3.340045e-08, -9.921479e-08, 1.032131e-08, 
    2.463878e-09, 1.852584e-09, 7.394959e-09, 3.725217e-09, 4.077498e-08, 
    1.526024e-08, 1.60957e-07, 4.47659e-08, -7.048067e-08, 2.195949e-07, 
    -2.212522e-08, -1.055692e-07, -7.256062e-10, 1.998177e-07, 2.674823e-07, 
    -3.838937e-08, -1.212128e-07, 5.066056e-09, 5.2801e-08, -1.716282e-07, 
    -1.534063e-07, -9.041556e-08, 6.793755e-09, 4.309805e-08, 5.306782e-08, 
    -2.091571e-08, 1.406357e-08, -5.973769e-08, 5.556281e-09, -5.250394e-08, 
    2.622158e-08, -1.854808e-07, -5.006922e-08, -5.013243e-08, -4.08665e-08, 
    -2.89387e-08, -3.270486e-09, 4.112678e-09, 3.251046e-09, -6.365042e-09, 
    2.014076e-10, 1.056776e-08, -3.171781e-09, -5.732446e-10, -1.36726e-08,
  2.830583e-07, 1.609766e-08, 1.202201e-07, 1.103113e-07, 1.329418e-07, 
    -1.257098e-08, 3.491039e-09, 4.036963e-09, 1.072062e-07, -7.080814e-09, 
    -4.757118e-08, 4.001339e-08, -7.910779e-08, 1.128074e-07, 2.70353e-09, 
    8.852862e-08, -2.235417e-07, 4.483957e-08, -3.128804e-09, -1.227382e-07, 
    2.176574e-08, -1.878759e-07, 9.405272e-08, -5.178339e-08, -1.834247e-07, 
    7.049169e-08, -4.553868e-08, -2.368114e-08, -1.025772e-07, -9.168815e-08, 
    -6.905515e-08, 3.485127e-09, -2.790779e-08, 9.777466e-09, 3.729127e-08, 
    5.925074e-09, -1.175476e-07, 1.141036e-08, -2.047312e-08, -9.13743e-08, 
    1.112621e-07, 2.06301e-07, 6.142369e-08, -6.079519e-08, -3.975458e-09, 
    -2.091366e-08, 5.055091e-08, -2.183012e-08, -1.411125e-08, 2.0732e-09, 
    6.293178e-09, -1.117853e-07, -7.463336e-08, 3.136339e-08, -3.920253e-08, 
    -1.559272e-09, 1.522324e-09, -2.192657e-07, -3.066248e-09, 7.16755e-08, 
    1.450814e-07, -1.394921e-07, 3.977491e-07, 1.391265e-07, -1.911491e-07, 
    -2.707583e-08, 2.499524e-08, -3.577276e-08, -3.302438e-08, -1.965265e-08, 
    -8.564808e-08, -1.309729e-07, -1.030876e-07, -2.632254e-08, 1.552532e-08, 
    4.30299e-09, 9.483117e-09, 3.575906e-09, -2.157694e-09, 2.357109e-08, 
    2.288391e-08, 1.572237e-07, 9.738301e-09, -8.200124e-08, 2.96605e-08, 
    -7.286246e-09, -1.702575e-07, 1.816096e-08, 1.739117e-07, 1.955066e-07, 
    -4.725081e-08, -1.114521e-07, 8.103541e-09, 1.226802e-07, -7.953753e-08, 
    3.546757e-08, -9.713284e-08, -7.696428e-09, 2.646715e-08, 4.241973e-08, 
    -1.457846e-08, 3.893049e-09, -1.579179e-07, 5.188276e-09, -2.579412e-08, 
    3.836527e-08, -1.649495e-07, -8.245917e-08, -8.851094e-08, -3.138751e-08, 
    -2.999121e-08, -5.135178e-09, 1.528349e-09, 4.069591e-09, -1.075415e-08, 
    1.200124e-09, 1.213336e-08, -2.877709e-09, -4.048744e-10, 1.649582e-07,
  1.340684e-07, 8.411405e-09, 2.003304e-07, 2.762676e-07, 6.610702e-08, 
    9.469164e-08, 1.704854e-08, 2.407906e-07, 7.888406e-08, 1.642101e-07, 
    9.334696e-08, 3.276801e-08, 2.535006e-07, 9.52902e-08, 1.267148e-08, 
    1.171338e-07, -2.292089e-07, 5.143437e-08, -7.484019e-09, -1.028209e-07, 
    6.105552e-10, -1.219789e-07, 1.388378e-07, -3.446138e-08, -2.878375e-08, 
    -1.215625e-08, -4.296049e-08, -1.421591e-08, -9.362094e-08, 
    -4.873442e-08, -6.777708e-08, 9.550263e-10, 1.645338e-08, -2.017958e-08, 
    -1.144377e-07, -8.348309e-09, -9.811898e-08, 9.208094e-09, -2.676614e-08, 
    -7.808592e-08, 1.165226e-07, 1.903359e-07, -6.144657e-08, -4.876079e-08, 
    -1.273003e-08, -5.665612e-08, 6.992536e-09, -1.063307e-07, -2.093901e-08, 
    1.983985e-09, 5.342869e-09, -1.59326e-07, -4.793502e-08, 2.858648e-08, 
    -3.161657e-08, -2.180855e-09, 4.426516e-08, -1.809224e-08, -4.338446e-09, 
    4.607686e-08, 3.162558e-08, -4.269606e-08, 3.717895e-08, 1.424238e-07, 
    -1.184877e-07, -2.528071e-08, 5.20771e-09, -3.694043e-08, -3.85217e-08, 
    -3.183624e-08, -7.80588e-08, -1.080129e-07, -1.998298e-07, -6.73578e-08, 
    1.440268e-08, 1.818591e-09, 1.906884e-09, -7.170598e-09, 4.557805e-09, 
    -6.254498e-08, 5.959123e-09, 1.414493e-07, 6.884125e-08, -7.86693e-08, 
    -2.209885e-08, 2.792711e-08, -1.975633e-07, 4.739724e-08, 1.481435e-07, 
    1.41515e-07, -5.716913e-09, -7.934874e-08, -1.121032e-08, 1.612137e-07, 
    -8.222685e-09, -3.498943e-08, -6.349843e-08, -4.314808e-08, 7.540791e-09, 
    1.129282e-08, -1.579753e-08, -1.701436e-07, -1.634068e-07, 3.504525e-09, 
    -8.020208e-09, 4.748466e-08, -1.651601e-07, -9.181548e-08, -9.911327e-08, 
    -2.921769e-08, -3.039264e-08, -6.007042e-09, 1.669491e-10, 4.162246e-09, 
    -1.14116e-08, 2.166985e-09, 4.922597e-09, -2.689518e-09, -2.278355e-10, 
    4.974498e-08,
  8.270956e-08, -6.33824e-07, 4.975118e-08, 2.023066e-07, 5.551431e-08, 
    7.600829e-08, 2.607396e-08, 8.147344e-08, -5.160427e-08, 9.850316e-08, 
    8.71953e-08, 4.11668e-08, 1.189353e-07, 5.543905e-08, 2.75013e-08, 
    1.137582e-07, -2.047925e-07, 3.621756e-08, 4.539771e-09, -1.806825e-08, 
    -4.504841e-09, -9.207952e-09, 3.206208e-08, -2.078775e-08, -3.293621e-09, 
    -3.296805e-08, -5.738252e-08, -1.711487e-08, -7.333767e-08, 2.46971e-08, 
    -4.367405e-08, 8.416418e-08, 1.375713e-08, -1.443141e-09, -2.017672e-07, 
    -1.224043e-08, -1.848322e-08, 6.511243e-09, -2.875652e-08, -2.835435e-08, 
    8.091344e-08, 5.946254e-08, -9.847204e-08, -4.131837e-08, -2.067827e-08, 
    -6.948608e-08, -2.718144e-08, -1.329579e-07, -2.030533e-08, 1.999865e-09, 
    4.494026e-09, -6.223456e-07, -2.34526e-08, 2.150493e-08, -2.660199e-08, 
    -1.793069e-09, 3.010415e-07, -4.545636e-08, -5.341228e-09, 3.943205e-08, 
    2.436764e-08, 1.096612e-08, 1.931983e-07, 1.543603e-07, -9.989165e-08, 
    -1.511353e-08, -6.963091e-09, -3.473701e-08, -2.704155e-08, 
    -2.968011e-08, -7.496999e-08, -5.870777e-08, -7.73972e-08, -6.072469e-09, 
    1.286795e-08, -2.870593e-09, -2.263971e-08, -1.128726e-08, 4.49343e-09, 
    4.818389e-08, -9.6191e-09, 1.130092e-07, 8.513274e-08, -4.679873e-08, 
    -8.576376e-08, 8.673589e-08, -3.015714e-07, 5.994809e-08, 1.21643e-07, 
    1.03706e-07, 4.82521e-09, -6.424074e-08, -7.696997e-09, 1.665513e-07, 
    2.716774e-09, -1.035076e-07, -3.548437e-08, -9.773657e-08, 1.425178e-09, 
    8.244108e-08, -1.064927e-08, -6.552814e-08, -1.353097e-07, 6.819342e-09, 
    -2.301647e-08, 5.809443e-08, -1.591668e-07, -9.456016e-08, -8.934796e-08, 
    -3.089701e-08, -3.016055e-08, -5.492439e-09, -6.025402e-10, 4.213462e-09, 
    -1.147873e-08, 4.473054e-09, 4.621256e-09, -2.442398e-09, -3.920135e-10, 
    1.140052e-08,
  6.203868e-08, -9.019993e-08, 3.795458e-08, -1.134595e-09, 1.153788e-07, 
    4.794106e-08, 5.35116e-08, -1.90438e-08, -2.933177e-08, 2.172339e-08, 
    1.820636e-07, 9.803432e-08, 3.854484e-08, -1.781859e-08, -2.300169e-08, 
    8.144783e-08, -1.707665e-07, -9.823339e-09, -3.020149e-08, 1.95161e-07, 
    -1.316141e-08, 1.05664e-08, 1.837975e-08, -1.493981e-08, 1.582657e-08, 
    -3.62154e-08, 3.438231e-09, -1.983165e-08, -4.383378e-08, 5.81507e-08, 
    8.973302e-09, 5.831987e-08, -4.841138e-08, 2.34229e-08, 8.91938e-08, 
    -5.645006e-09, 2.017902e-08, 4.969777e-09, 1.414048e-08, -2.128878e-08, 
    7.505628e-08, 3.44445e-08, -7.794671e-08, -2.165803e-08, -1.124624e-08, 
    -7.616154e-08, -4.798807e-08, -1.210103e-07, -2.005561e-08, 1.979529e-09, 
    3.791001e-09, -1.098387e-07, -8.592486e-09, 2.517777e-08, -2.249869e-08, 
    -1.237538e-09, 1.477293e-07, 5.989746e-08, -6.178993e-09, -3.656311e-08, 
    2.032539e-08, 3.196703e-08, 2.376748e-08, 1.19663e-07, -1.419414e-07, 
    -2.517834e-08, 3.706418e-09, -5.76199e-09, 1.214312e-08, -3.697085e-08, 
    -6.514153e-08, 1.225201e-07, 2.128945e-08, 1.560886e-08, 1.22191e-08, 
    -9.624614e-09, 4.786826e-08, -1.971134e-08, 1.039587e-08, 6.375501e-08, 
    -1.096873e-08, 9.271536e-08, 3.115036e-08, -4.277922e-09, -2.119884e-08, 
    2.985496e-08, -1.416269e-07, -4.451044e-08, 9.874358e-08, 7.938098e-08, 
    5.275979e-09, -6.691589e-08, -5.582706e-09, 1.68154e-07, -4.689559e-08, 
    -1.272557e-07, -1.020897e-07, -9.203654e-08, 1.380329e-08, 8.756588e-08, 
    6.028733e-08, -9.031282e-10, -2.580337e-08, 7.43853e-09, -4.987373e-08, 
    5.241145e-08, -1.352994e-07, -9.621397e-08, -8.924997e-08, -3.211028e-08, 
    -2.815398e-08, -5.722654e-09, -1.006697e-09, 4.178901e-09, -1.16388e-08, 
    7.692393e-09, 2.110767e-09, -2.226159e-09, -7.052279e-10, -5.167669e-08,
  5.58145e-08, -7.115403e-08, 3.343627e-08, -1.000348e-08, 1.227653e-08, 
    -6.818198e-09, 1.345085e-07, -3.022564e-08, -3.351187e-08, -2.961525e-08, 
    -2.600217e-08, 1.148902e-08, -7.872529e-09, -2.376379e-08, -3.060183e-08, 
    5.602892e-08, -1.426769e-07, -2.700313e-08, 4.412865e-08, -3.925282e-08, 
    -1.230109e-08, 1.634368e-08, 9.850112e-09, -1.165103e-08, 2.549365e-08, 
    -3.727854e-08, -4.981558e-08, -2.46078e-08, 2.195014e-08, 8.107617e-08, 
    7.171877e-09, 8.478258e-08, 5.889268e-08, 1.52732e-08, 7.956686e-08, 
    4.685091e-09, 3.082144e-08, 5.268888e-09, -1.736736e-07, -2.681903e-08, 
    4.225009e-08, 1.998086e-08, -6.772143e-08, -4.850643e-09, -1.346604e-08, 
    -8.369165e-08, -6.09262e-08, -1.111642e-07, -1.896113e-08, 1.895621e-09, 
    3.294957e-09, -3.200836e-08, 2.793115e-09, 2.986464e-08, -1.811202e-08, 
    3.821015e-10, 1.464583e-07, 4.409281e-08, -7.002143e-09, -4.714066e-08, 
    1.774362e-08, 3.900567e-08, -3.609244e-08, 8.887584e-08, -9.159285e-08, 
    -6.689191e-08, 3.643663e-11, 3.497638e-08, 3.433968e-09, -5.404564e-08, 
    -7.758257e-08, 3.008035e-07, -6.552324e-08, 1.19374e-08, 1.209502e-08, 
    -2.019573e-08, -1.257669e-08, -1.049742e-08, 1.730074e-08, 1.412517e-07, 
    4.236938e-09, 7.271056e-08, 1.321723e-08, 6.568882e-09, 7.370488e-09, 
    -6.609156e-08, -6.859722e-08, -9.635772e-08, 9.786504e-08, 6.509754e-08, 
    5.19077e-09, -7.449586e-08, -9.838772e-09, 1.55892e-07, -6.725145e-10, 
    -1.426998e-07, -1.724039e-07, -1.140065e-07, 9.447433e-09, 5.148426e-08, 
    2.014921e-07, 1.208073e-08, 2.231599e-08, 7.118629e-09, -3.523411e-08, 
    9.101825e-09, -1.388664e-07, -9.358968e-08, -8.618525e-08, -3.254337e-08, 
    -2.797043e-08, -5.818322e-09, -9.186465e-10, 4.108358e-09, -1.036659e-08, 
    1.293724e-08, 2.217888e-10, -2.583118e-09, -8.424124e-10, -6.353895e-08,
  5.318202e-08, -6.744233e-08, 3.269543e-08, -1.257661e-08, 6.121695e-09, 
    -1.355363e-08, 1.270996e-08, -4.443211e-08, -3.956143e-08, -4.173739e-08, 
    -6.406731e-08, -6.583844e-08, -1.990099e-08, -2.707418e-08, 
    -3.271725e-08, 4.666978e-08, -8.760715e-08, 4.332549e-09, 8.004555e-08, 
    -6.186599e-08, -1.217529e-08, 2.099728e-08, 6.165806e-09, -9.653718e-09, 
    2.366426e-08, -3.774176e-08, -5.752815e-08, -9.222458e-08, 2.13472e-08, 
    -2.965487e-08, 1.009289e-08, 6.729806e-09, 6.662322e-08, 1.452941e-08, 
    5.08328e-08, 2.826039e-08, 2.901875e-08, 5.686601e-09, -1.764861e-07, 
    -1.928824e-08, 1.453091e-08, 9.455789e-09, -6.146672e-08, -4.319626e-09, 
    -1.314891e-08, -9.075063e-08, -6.841515e-08, -1.045106e-07, 
    -1.939432e-08, 2.237115e-09, 2.926654e-09, -6.606001e-09, 1.211771e-08, 
    3.44284e-08, -1.400434e-08, -9.566179e-10, 2.004115e-07, 4.252094e-08, 
    -7.61537e-09, -2.6816e-08, 1.605156e-08, 4.154936e-08, -4.251649e-08, 
    4.422193e-08, -4.512135e-08, -7.989343e-09, 2.468971e-08, 4.152821e-08, 
    3.835112e-09, -5.487072e-08, -7.82187e-08, 1.891967e-07, -8.318182e-08, 
    1.403464e-08, 1.128258e-08, -2.35832e-08, -2.035887e-08, -5.937835e-09, 
    1.924672e-08, 2.066652e-07, -9.429357e-09, 5.857889e-08, 9.099438e-09, 
    7.940457e-09, 1.326748e-08, -4.078493e-08, -4.986703e-08, -4.163201e-08, 
    1.019074e-07, 5.827297e-08, 5.191396e-09, -6.567534e-08, -1.780066e-08, 
    1.38254e-07, 1.490434e-08, -1.487929e-07, -1.982591e-07, -8.725351e-08, 
    1.168826e-08, 1.859737e-08, 1.120636e-07, 1.875701e-08, 4.023153e-08, 
    6.589616e-09, 3.314437e-08, 4.520189e-09, -2.176328e-07, -7.812503e-08, 
    -7.871336e-08, -3.112439e-08, -2.818956e-08, -3.168452e-09, 
    -1.152102e-09, 4.067374e-09, -8.746611e-09, 6.852964e-09, 1.068003e-09, 
    -1.901984e-09, -4.233982e-10, -6.848711e-08,
  5.204873e-08, -6.491933e-08, 3.188137e-08, -1.148209e-08, 2.739455e-09, 
    -1.636243e-08, -1.592053e-08, -4.947577e-08, -4.148711e-08, 
    -4.696705e-08, -8.467742e-08, -8.268461e-08, -2.428811e-08, 
    -2.796929e-08, -3.346821e-08, 4.294927e-08, -2.982747e-08, 1.398291e-09, 
    9.242022e-08, -7.320347e-08, -1.213851e-08, 2.51726e-08, 4.860397e-09, 
    -8.696759e-09, 2.426333e-08, -3.786005e-08, -4.519092e-08, 9.820781e-09, 
    2.142275e-08, -4.880479e-08, 8.472682e-09, -1.762936e-08, 9.603679e-08, 
    2.528458e-08, 5.294663e-08, 6.108172e-08, 2.47698e-08, 5.838132e-09, 
    -1.729337e-07, -1.306735e-08, 5.161951e-09, 2.73684e-09, -6.017183e-08, 
    -7.376391e-09, -3.640019e-08, -9.191166e-08, -7.227686e-08, -9.53342e-08, 
    -2.017297e-08, 4.363599e-09, 2.682583e-09, 2.226386e-09, 1.785113e-08, 
    3.73164e-08, -1.095262e-08, -1.438877e-09, 2.188089e-07, 4.1032e-08, 
    -8.173302e-09, -1.528591e-09, 1.497102e-08, 4.3645e-08, -4.789757e-08, 
    3.047729e-08, -2.233588e-08, -6.00831e-08, -3.457859e-08, 2.310759e-08, 
    -8.691188e-09, -4.774853e-08, -5.00275e-08, -5.099395e-08, -7.570253e-08, 
    1.411632e-08, 1.054601e-08, -2.114956e-08, -2.152399e-08, -8.799361e-11, 
    1.770317e-08, 2.199803e-07, -1.163289e-08, 4.993352e-08, 7.908909e-09, 
    7.936762e-09, 2.194741e-08, -4.461697e-09, -5.790315e-08, -1.879113e-08, 
    1.007784e-07, 5.571906e-08, 5.273762e-09, -7.230263e-08, -2.02254e-08, 
    1.206625e-07, 4.725877e-08, -1.516965e-07, -2.093022e-07, -8.937775e-09, 
    1.557856e-08, -1.732573e-08, 8.974411e-08, 2.221812e-08, 6.643209e-08, 
    5.14482e-09, 4.656596e-08, 2.508199e-08, -2.359316e-07, -5.60006e-08, 
    -6.626868e-08, -2.833787e-08, -2.824851e-08, -1.414207e-09, 
    -1.295632e-09, 4.072092e-09, -4.031733e-09, -1.174953e-10, 2.858286e-09, 
    -1.49673e-09, -1.036256e-10, -7.071452e-08,
  5.166578e-08, -6.31378e-08, 4.15896e-08, -1.462479e-08, 1.676881e-09, 
    -1.814044e-08, -1.827607e-08, -5.157733e-08, -4.171784e-08, 
    -4.865058e-08, -9.270502e-08, -9.024791e-08, -2.617605e-08, 
    -3.085097e-08, -3.375055e-08, 2.354756e-08, 8.625189e-10, -6.581331e-10, 
    9.235396e-08, -7.809638e-08, -1.221429e-08, 2.824936e-08, 3.724153e-09, 
    -8.570964e-09, 2.34113e-08, -3.780019e-08, -4.889637e-08, 2.470631e-08, 
    2.010131e-08, -8.318921e-09, 1.332216e-08, 4.298397e-08, 9.227267e-08, 
    2.979107e-08, 5.072434e-08, 7.42325e-08, 2.031733e-08, 5.125671e-09, 
    8.174266e-08, -7.815618e-09, -3.313454e-08, -9.073347e-10, -6.016302e-08, 
    -6.217711e-09, -4.411629e-08, -9.942312e-08, -7.445925e-08, 
    -9.044905e-08, -1.907056e-08, -2.286008e-09, 2.531479e-09, 5.513243e-09, 
    2.150006e-08, 3.878063e-08, -8.770383e-09, -2.775323e-09, 2.276663e-07, 
    3.925457e-08, -8.804193e-09, 2.231289e-08, 1.444209e-08, 4.46305e-08, 
    -5.033337e-08, 2.041209e-08, -9.578412e-09, 7.777658e-09, -9.60631e-09, 
    -4.590333e-09, -1.20906e-08, -6.720302e-08, -5.279878e-08, -1.226341e-07, 
    -1.037499e-07, 1.359604e-08, 9.771647e-09, -1.621072e-08, -2.208091e-08, 
    2.109687e-09, 1.512601e-08, 2.301825e-07, -1.320404e-08, 4.436335e-08, 
    7.399649e-09, 7.728204e-09, 2.862589e-08, -6.902951e-09, -5.961931e-08, 
    -1.08821e-08, 1.048028e-07, 5.603562e-08, 5.641937e-09, -4.769911e-08, 
    -2.631958e-08, 1.133814e-07, 5.228537e-08, -1.522977e-07, -2.132674e-07, 
    -1.848025e-08, 1.760577e-08, -3.016651e-08, 8.370159e-08, 2.758895e-08, 
    7.099766e-08, 4.647646e-09, 5.204333e-08, 4.515516e-08, -1.882275e-07, 
    -2.787783e-08, -4.711842e-08, -2.307809e-08, -2.273305e-08, 
    -4.952199e-10, -1.135959e-09, 4.024969e-09, 1.069793e-09, 6.566552e-10, 
    2.783054e-10, -1.200629e-09, -2.27125e-10, -7.12148e-08,
  4.971145e-08, -6.160775e-08, 4.542807e-08, -1.223663e-08, 1.936485e-09, 
    -1.915004e-08, -2.09829e-08, -5.220494e-08, -4.13275e-08, -4.781617e-08, 
    -9.592583e-08, -9.398758e-08, -2.701398e-08, -3.064639e-08, -3.40188e-08, 
    -9.863385e-09, 1.193719e-08, -2.08081e-09, 9.385892e-08, -8.062631e-08, 
    -1.228392e-08, 2.855546e-08, 2.67238e-09, -8.610357e-09, 2.249243e-08, 
    -3.78414e-08, -4.0168e-08, -1.207663e-07, 1.962593e-08, -5.851751e-08, 
    1.768746e-08, 6.555257e-08, 1.094132e-07, 2.965129e-08, 4.907525e-08, 
    6.957504e-08, 1.654896e-08, 1.427821e-09, 2.032535e-07, -7.209849e-09, 
    -7.403918e-08, -2.182958e-09, -6.029214e-08, -1.029404e-09, 
    -9.430266e-09, -1.070492e-07, -7.562204e-08, -8.777826e-08, 
    -1.655691e-08, -6.401137e-10, 2.467445e-09, 6.963603e-09, 2.375898e-08, 
    3.888257e-08, -7.193273e-09, -5.281834e-09, 2.36372e-07, 3.876281e-08, 
    -9.558647e-09, 3.905882e-08, 1.413201e-08, 4.505199e-08, -5.175383e-08, 
    1.357692e-08, -4.654601e-09, 2.02935e-08, -4.864154e-08, 3.923566e-08, 
    -1.542759e-08, -7.135185e-08, -4.087309e-08, -1.448448e-07, 
    -1.181846e-07, 1.290113e-08, 9.023498e-09, 6.221683e-09, -2.248026e-08, 
    3.246441e-09, 1.312636e-08, 2.3447e-07, -7.600704e-09, 4.073629e-08, 
    7.163408e-09, 7.525671e-09, 3.253371e-08, 3.757975e-09, -5.986811e-08, 
    -6.814332e-09, 1.204929e-07, 5.904809e-08, 5.618801e-09, -3.865692e-08, 
    -2.046508e-08, 1.075391e-07, 6.254282e-08, -1.521084e-07, -2.111994e-07, 
    -1.498864e-08, 1.835912e-08, -3.788908e-08, 7.887826e-08, 3.040438e-08, 
    6.875267e-08, 4.659618e-09, 5.401847e-08, 4.651787e-08, -8.223213e-08, 
    2.448303e-09, -2.522967e-08, -1.582515e-08, -1.958523e-08, 1.8685e-09, 
    -4.473577e-11, 4.04151e-09, 2.905551e-09, -7.316316e-10, -1.925613e-09, 
    -1.795719e-10, -5.929337e-10, -7.04967e-08,
  4.953881e-08, -6.156415e-08, 9.16516e-08, -1.083731e-08, 2.284196e-09, 
    -1.994999e-08, -2.523655e-08, -5.273307e-08, -3.82571e-08, -4.447838e-08, 
    -9.679241e-08, -9.550024e-08, -2.712466e-08, -3.065554e-08, 
    -3.373407e-08, -4.321919e-08, 1.521991e-08, -2.597744e-09, 9.369644e-08, 
    -8.184008e-08, -1.203557e-08, 2.991862e-08, 1.776016e-09, -9.539463e-09, 
    2.101706e-08, -3.777416e-08, -3.404261e-08, -1.10981e-07, 1.949923e-08, 
    -7.050983e-08, 2.126558e-08, 7.07455e-08, 1.211512e-07, 1.833746e-08, 
    4.661081e-08, 5.778372e-08, 1.432937e-08, 1.759119e-09, -3.860885e-08, 
    -6.517974e-09, -1.363479e-07, -1.703029e-09, -5.969613e-08, 2.764859e-09, 
    4.529284e-10, -1.121695e-07, -7.616592e-08, -8.742407e-08, -1.325582e-08, 
    -5.16799e-10, 2.3757e-09, 7.711947e-09, 2.494239e-08, 4.103222e-08, 
    -5.805569e-09, -7.793176e-09, 2.391608e-07, 3.699733e-08, -1.050395e-08, 
    5.370295e-08, 1.397075e-08, 4.565186e-08, -5.217305e-08, 8.284147e-10, 
    -6.595542e-09, 1.87872e-08, -5.000493e-08, 4.020137e-08, -1.758337e-08, 
    -6.878759e-08, -2.448883e-08, -1.542659e-07, -1.275282e-07, 1.144031e-08, 
    8.293419e-09, 1.912292e-08, -2.221741e-08, 3.98137e-09, 1.224159e-08, 
    2.350038e-07, -3.084892e-09, 3.877684e-08, 7.195013e-09, 7.339736e-09, 
    2.986405e-08, 7.729341e-09, -5.920333e-08, -4.291792e-09, 1.193493e-07, 
    6.358277e-08, 6.038476e-09, -3.552802e-08, -1.927575e-08, 1.05187e-07, 
    6.86606e-08, -1.520428e-07, -2.092268e-07, -5.886363e-09, 1.992544e-08, 
    -3.951798e-08, 7.798428e-08, 3.157017e-08, 6.624281e-08, 4.75098e-09, 
    5.451273e-08, 4.700564e-08, 7.122298e-08, 3.576804e-08, -4.597723e-09, 
    -8.190568e-09, -1.56823e-08, 4.588401e-09, 1.697458e-09, 4.021786e-09, 
    4.779281e-09, 8.1194e-10, -2.209347e-09, -1.275851e-10, -3.176552e-10, 
    -6.805465e-08,
  4.927165e-08, -5.960658e-08, 1.133944e-07, -8.524921e-09, 3.813784e-08, 
    -2.115917e-08, -2.78294e-08, -5.198376e-08, -3.633977e-08, -4.473532e-08, 
    -9.600592e-08, -9.50389e-08, -2.651268e-08, -2.883621e-08, -3.309367e-08, 
    -4.052785e-08, 1.580326e-08, -4.144397e-09, 9.41847e-08, -8.196059e-08, 
    -1.180933e-08, 3.050855e-08, 8.742518e-10, -1.149613e-08, 1.891567e-08, 
    -3.767241e-08, -3.467369e-08, -1.092619e-07, 1.976764e-08, -8.375082e-08, 
    2.453135e-08, 7.019548e-08, 1.280229e-07, -4.436515e-09, 4.593551e-08, 
    4.379626e-08, 9.895814e-09, 9.758594e-11, -1.751354e-07, -6.690652e-09, 
    -2.316239e-07, 1.955414e-10, -5.892312e-08, 5.360846e-09, -1.296939e-09, 
    -1.185953e-07, -7.636362e-08, -8.911528e-08, -1.378692e-08, -1.54467e-09, 
    2.390109e-09, 8.092115e-09, 2.580125e-08, 4.504848e-08, -3.825323e-09, 
    -6.672508e-09, 2.410353e-07, 3.572142e-08, -1.179399e-08, 6.334569e-08, 
    1.395028e-08, 4.62984e-08, -5.089453e-08, -1.374207e-08, -9.43628e-09, 
    2.154934e-08, -4.577248e-08, 6.317214e-08, -1.521823e-08, -6.362347e-08, 
    -9.202267e-09, -1.556436e-07, -1.290761e-07, 1.082549e-08, 7.297057e-09, 
    3.378773e-10, -2.191409e-08, 3.917165e-09, 1.147435e-08, 2.318767e-07, 
    -4.401159e-09, 3.769521e-08, 9.558278e-09, 7.113954e-09, 2.349827e-08, 
    1.138051e-08, -5.799484e-08, -2.31546e-09, 1.208727e-07, 6.941565e-08, 
    5.793709e-09, -3.199695e-08, -1.878263e-08, 8.979694e-08, 7.360006e-08, 
    -1.511156e-07, -2.061886e-07, -2.623324e-09, 1.983608e-08, -4.013841e-08, 
    7.894607e-08, 3.079718e-08, 7.333433e-08, 4.848872e-09, 5.363984e-08, 
    4.506012e-08, 1.077735e-07, 6.491621e-08, 1.203307e-08, -1.518174e-09, 
    -1.129081e-08, 8.569941e-09, 3.888317e-09, 6.096911e-09, 6.133632e-09, 
    -2.525053e-09, 2.230095e-09, -2.354835e-09, -8.645173e-10, -6.433288e-08,
  4.903131e-08, -5.426557e-08, 1.181533e-07, -3.158107e-09, 4.43265e-08, 
    -2.268166e-08, -2.99317e-08, -4.964249e-08, -3.397508e-08, -4.236017e-08, 
    -9.23161e-08, -9.059738e-08, -2.437855e-08, -2.391744e-08, -3.115929e-08, 
    -3.753848e-08, 1.653066e-08, -5.697018e-09, 8.856496e-08, -8.018446e-08, 
    -1.196838e-08, 2.871855e-08, -1.250555e-10, -1.224146e-08, 1.497472e-08, 
    -3.740263e-08, -3.113848e-08, -1.105076e-07, 2.083425e-08, -7.716335e-08, 
    2.856098e-08, 6.699406e-08, 1.2481e-07, -2.961281e-08, 4.514334e-08, 
    3.687114e-08, 1.003326e-08, 1.151506e-10, -1.941655e-07, -7.826168e-09, 
    -4.169185e-07, 4.429808e-09, -5.721319e-08, 3.506962e-09, -4.551111e-09, 
    -1.24125e-07, -7.634623e-08, -9.32755e-08, -1.557751e-08, -4.878856e-09, 
    2.493636e-09, 8.19125e-09, 2.672741e-08, 4.805306e-08, -9.772663e-10, 
    -6.927905e-09, 2.26394e-07, 2.702107e-08, -1.384205e-08, 6.70499e-08, 
    1.405158e-08, 4.723631e-08, -4.662581e-08, -3.294797e-08, -1.856104e-08, 
    2.134345e-08, -4.706703e-08, 6.689345e-08, -7.551648e-09, -6.435187e-08, 
    5.949914e-09, -1.97202e-07, -1.19271e-07, 7.628273e-09, 5.626724e-09, 
    -5.703782e-09, -2.130243e-08, 3.744844e-09, 6.495796e-09, 2.200401e-07, 
    -6.628454e-09, 3.774873e-08, 1.100625e-08, 6.94456e-09, 2.127945e-08, 
    4.733351e-09, -5.587049e-08, -2.116849e-10, 1.185574e-07, 8.089455e-08, 
    5.479706e-09, -2.843124e-08, -1.75956e-08, 7.818786e-08, 7.089238e-08, 
    -1.479027e-07, -1.984434e-07, 3.508603e-09, 1.842375e-08, -3.858317e-08, 
    7.780375e-08, 2.711734e-08, 7.04819e-08, 4.86498e-09, 4.980211e-08, 
    3.871833e-08, 1.110088e-07, 7.940014e-08, 1.496778e-08, 1.19519e-09, 
    -7.229119e-09, 1.436513e-08, 9.832434e-09, 1.131627e-08, 7.283347e-09, 
    -3.257696e-10, 4.023534e-08, 1.375994e-09, -5.862887e-09, -5.733818e-08,
  3.446799e-13, 4.300897e-14, -1.753807e-13, -3.633421e-13, -3.538563e-13, 
    -1.570426e-13, 2.545201e-13, 1.065312e-13, -2.767669e-13, -2.00539e-13, 
    -4.697948e-13, -5.748564e-13, 2.39716e-13, 1.773635e-14, -1.040004e-13, 
    1.387841e-13, -7.51801e-13, -1.308467e-13, -1.315635e-13, -1.284254e-13, 
    -1.94583e-12, -2.475496e-12, -6.430807e-14, 5.739497e-13, -1.282557e-12, 
    -1.900151e-13, 1.609106e-13, 9.396559e-14, 6.188501e-14, 7.188945e-14, 
    -3.050115e-14, 3.067236e-14, 3.775378e-14, 2.014006e-13, 4.128115e-14, 
    3.612441e-13, -5.59297e-13, -3.368272e-12, 2.72692e-14, 3.213058e-12, 
    2.298948e-13, -7.20349e-14, -1.705905e-13, 2.65163e-13, 1.137971e-13, 
    4.721511e-13, 5.338034e-13, 1.587444e-12, 8.619935e-13, 1.340315e-12, 
    -5.139416e-13, -3.523681e-14, 1.990189e-12, -6.518992e-13, 5.021289e-14, 
    -4.989662e-13, 2.880441e-13, 2.023415e-13, 1.276777e-13, 3.705946e-13, 
    9.474537e-13, -1.610186e-13, 5.380253e-13, -1.914522e-12, -3.802779e-13, 
    3.329098e-13, -8.124365e-14, -3.301351e-13, -1.125156e-14, 8.227237e-14, 
    -1.345926e-13, -7.472412e-14, 7.560632e-14, 3.384418e-13, -1.247063e-12, 
    -6.071229e-13, -1.538443e-13, -9.914854e-13, -1.400826e-12, 
    -1.547843e-13, 4.857807e-14, 1.350339e-12, -4.313481e-13, -5.958526e-13, 
    3.193387e-14, 8.412611e-14, -3.455108e-13, 8.105178e-13, 1.661521e-12, 
    6.491071e-13, 3.131953e-13, 2.057114e-12, -7.770231e-13, -9.624789e-14, 
    -2.16057e-13, -4.0491e-13, 3.004785e-13, -7.872333e-14, 1.89724e-13, 
    -3.556957e-13, -5.763276e-13, 4.06125e-13, -9.685324e-13, 2.17412e-13, 
    9.234387e-15, 3.733669e-13, 5.788955e-15, -5.279393e-13, -6.430571e-13, 
    -1.984821e-13, 9.166984e-15, -7.987311e-14, -2.126898e-14, -9.929794e-15, 
    4.531738e-13, -3.613456e-12, -3.71223e-13, -6.61266e-13, 1.933037e-12, 
    6.675825e-14,
  3.70461e-13, 2.683964e-13, 1.770327e-13, 1.275379e-13, 8.761511e-14, 
    5.374604e-14, -4.98479e-14, -3.108878e-13, -1.136497e-13, -2.95671e-13, 
    -3.493155e-13, -1.63712e-13, -2.710435e-13, -4.394112e-13, -3.867215e-13, 
    3.171501e-13, 8.174496e-14, -2.489214e-13, -2.795625e-13, -3.805238e-14, 
    7.76688e-14, -3.861904e-13, -2.465668e-14, -1.294626e-13, -2.665974e-13, 
    -5.181435e-13, -6.789085e-13, 5.960301e-14, 8.727922e-14, 2.774094e-13, 
    9.294207e-14, -5.680436e-14, -1.483338e-13, -3.184754e-13, -8.944232e-14, 
    8.842967e-14, -5.35406e-13, -2.645126e-13, -1.541546e-15, -1.298683e-12, 
    -9.091551e-13, 1.039657e-13, -2.638347e-13, 2.151754e-13, -8.903726e-13, 
    -7.290542e-13, -1.058995e-12, 9.547694e-13, -6.700765e-15, 4.324396e-13, 
    -1.538602e-13, -1.374566e-13, 1.159862e-12, 1.369083e-12, 1.047405e-12, 
    -4.774958e-13, 6.319194e-14, -1.341717e-12, -2.530677e-13, 5.622747e-15, 
    4.537888e-14, 2.145897e-13, -1.460639e-13, -6.752341e-14, -9.513707e-14, 
    -1.251455e-13, 5.397915e-14, -1.253938e-13, -2.743941e-13, -3.459612e-13, 
    -1.119581e-12, 2.290802e-13, -5.173017e-13, -8.564723e-14, 1.324539e-13, 
    -5.296943e-13, 3.246323e-13, 1.380296e-12, -7.193178e-12, -1.322299e-13, 
    2.382339e-14, -1.817542e-13, -2.658812e-13, -1.302428e-13, -2.912002e-13, 
    5.917587e-13, -3.033076e-13, 1.484303e-13, -1.144643e-12, -1.950481e-13, 
    4.183061e-14, -1.382662e-13, 1.452668e-13, -5.807905e-13, 1.175756e-13, 
    2.369878e-13, 6.257669e-14, -1.186977e-13, 4.039507e-14, 1.155898e-12, 
    -8.712679e-13, 7.203452e-13, -2.71387e-13, -4.599547e-12, 1.263024e-13, 
    4.32073e-13, 8.034153e-13, 1.888171e-12, 1.390496e-12, 8.105602e-13, 
    4.250065e-13, 2.53079e-13, 1.022743e-13, 6.518476e-14, 4.450365e-13, 
    2.22772e-12, -9.70191e-13, -2.020404e-12, -4.847072e-14, 2.699439e-13,
  -2.607636e-14, -3.014256e-14, -8.305856e-14, -1.821043e-13, -2.701311e-13, 
    -2.627343e-13, -5.838385e-14, 2.980255e-13, 3.759076e-13, 1.664918e-13, 
    1.820766e-14, -2.506606e-13, -2.482181e-13, 1.157685e-13, 5.1259e-13, 
    6.094916e-13, 2.307293e-13, 4.503203e-13, 2.509104e-14, -8.580359e-13, 
    -5.862255e-13, -6.286083e-13, -7.220613e-13, -5.092593e-13, 
    -3.669981e-13, -3.165662e-13, 2.583073e-13, -1.379452e-14, -1.066924e-13, 
    5.294376e-14, 2.889355e-14, 2.781109e-14, -1.736111e-14, -7.024936e-14, 
    6.68493e-14, 1.309647e-13, -5.177289e-13, -8.057686e-13, 1.936923e-13, 
    -1.75438e-12, 6.220968e-13, 6.330075e-13, 1.331574e-13, 3.394268e-13, 
    2.519235e-13, 4.622275e-13, -1.887782e-12, -8.743319e-13, 2.554623e-13, 
    1.952397e-13, -1.649497e-13, -4.210798e-13, -5.983728e-13, -2.400975e-11, 
    2.951316e-13, 1.007548e-12, 3.831657e-13, -2.046226e-12, -1.242952e-12, 
    2.315212e-12, 8.308909e-13, -5.055678e-14, 2.888939e-13, 2.922523e-13, 
    4.009654e-13, 7.306655e-14, -8.160139e-15, -1.286748e-13, 3.871903e-15, 
    4.52971e-14, -1.39784e-12, 1.737777e-13, 9.652557e-13, -6.421252e-14, 
    -2.940315e-13, -2.349287e-12, -1.098472e-12, 2.220377e-13, -2.270685e-12, 
    -6.064871e-13, 3.632442e-13, 1.340145e-12, -2.916278e-13, -3.756856e-13, 
    -1.365991e-13, -4.805184e-13, -2.535624e-12, -2.667727e-13, 
    -2.130521e-12, -1.941697e-12, -1.127431e-13, -6.752821e-13, 2.69073e-13, 
    -2.552453e-12, 1.346145e-14, 2.374975e-13, 3.078371e-13, -1.83159e-13, 
    7.979312e-13, 1.517558e-12, 8.370943e-13, 1.33114e-13, 3.304631e-13, 
    -1.010451e-12, 2.464834e-13, 4.045514e-13, 3.91645e-13, -2.418898e-14, 
    -2.666201e-13, -6.39877e-13, -6.757234e-13, -1.044442e-13, 2.112199e-14, 
    1.776357e-13, 1.418449e-13, 3.337036e-12, 1.155469e-11, 3.91911e-12, 
    -4.484841e-13, -7.234907e-13,
  1.797174e-14, -2.692291e-14, -9.532652e-14, -8.149037e-14, -3.458345e-14, 
    4.10505e-14, 1.284806e-13, 2.58113e-13, 2.989414e-13, 3.860939e-13, 
    9.686696e-15, 5.330181e-13, 1.356831e-13, 1.088712e-13, -7.785439e-15, 
    3.689146e-13, 4.469245e-13, 3.930814e-13, 3.82026e-13, 4.399814e-13, 
    -8.720802e-14, -4.623663e-13, -7.056439e-13, 8.493206e-15, 1.372472e-12, 
    1.353473e-12, -1.422473e-14, -3.185091e-13, -4.08118e-13, -3.309297e-13, 
    1.011274e-13, 6.661338e-14, 6.189216e-13, 2.669254e-13, -4.194561e-13, 
    -2.14842e-13, -1.630283e-12, 1.416865e-12, -6.814826e-13, -4.584333e-13, 
    3.399753e-13, 3.865797e-13, 5.330458e-13, 3.72497e-13, 3.365364e-14, 
    -9.413165e-13, -2.435378e-12, -7.418545e-13, 8.876372e-13, -2.132921e-13, 
    -1.032273e-12, 1.931705e-12, -4.682144e-13, -1.766087e-14, 2.973413e-13, 
    1.366532e-12, -3.299139e-12, -9.613727e-13, 1.270511e-13, 1.911084e-12, 
    -1.969258e-14, -4.067718e-13, 1.173922e-12, 5.286966e-13, 5.012352e-13, 
    7.082529e-13, 4.480305e-13, 5.900697e-13, 6.778467e-13, -7.760459e-14, 
    -6.482315e-14, 6.201567e-13, 9.508366e-13, -2.028516e-13, -4.738876e-13, 
    -2.013389e-12, 1.770702e-13, 2.582722e-12, -8.240595e-12, -7.134571e-14, 
    1.225325e-12, -5.748478e-13, -7.564088e-14, 9.231782e-13, 1.07081e-13, 
    -1.428441e-13, -3.306105e-13, 3.354539e-13, -1.081844e-12, -1.047988e-12, 
    -3.466116e-13, -3.535738e-12, -2.174511e-13, 9.069245e-13, 4.654888e-13, 
    -3.263893e-11, 1.809414e-12, 1.205702e-13, -5.285106e-12, -1.871281e-13, 
    -1.054851e-12, -5.933275e-14, 2.964295e-13, -1.178866e-13, -1.013079e-15, 
    -1.94289e-16, 4.349299e-14, -7.05172e-13, -3.152895e-13, 1.011552e-13, 
    -3.83138e-13, -2.572526e-13, -2.250422e-13, -9.282852e-14, 1.475209e-14, 
    1.902194e-12, -7.607179e-13, 1.168025e-12, -1.107673e-13, 1.64771e-13,
  -1.826456e-13, 4.926476e-13, 4.859585e-13, 4.278383e-13, 3.345241e-13, 
    9.924006e-14, -2.136763e-13, 2.219197e-13, 9.169054e-14, -6.117468e-13, 
    3.113759e-13, 3.098494e-13, 4.361789e-14, -4.552331e-13, 2.865763e-14, 
    2.721851e-13, 4.863138e-13, 9.747064e-13, 7.002003e-13, 7.445017e-13, 
    7.07337e-13, 6.632195e-14, 8.733292e-14, 5.751927e-13, 7.351481e-13, 
    2.705752e-13, 3.722161e-13, 2.204487e-13, 2.844947e-15, 9.743595e-14, 
    6.991213e-13, -1.0872e-12, -5.438289e-13, 5.285355e-13, -6.471074e-13, 
    6.204759e-14, -1.114681e-12, -9.788004e-14, -1.554992e-12, -6.086825e-13, 
    -1.183356e-12, -3.80182e-13, 6.334794e-13, 1.825389e-13, -1.218678e-12, 
    -4.411332e-13, -1.861844e-13, 2.446376e-13, -5.886097e-13, 1.420478e-11, 
    -3.386354e-13, 9.738738e-13, 2.133016e-14, -1.347092e-12, 3.677267e-14, 
    1.076708e-12, -5.202991e-12, -2.217429e-12, -2.814304e-13, 7.208366e-13, 
    7.748663e-13, -7.445849e-13, -8.181372e-13, 5.095341e-13, 5.999951e-13, 
    -3.842343e-13, 1.807027e-13, 2.014361e-13, 1.618844e-13, 1.143544e-12, 
    9.767326e-13, -7.942258e-14, 3.769346e-13, -3.549244e-13, -5.531353e-13, 
    -1.020087e-12, -5.878804e-13, -4.488077e-13, -2.740484e-12, 
    -5.821732e-14, 4.434647e-13, 1.215748e-12, 3.933937e-13, 1.229641e-12, 
    5.236089e-14, -2.405756e-12, -4.314604e-14, 5.947881e-13, -1.085606e-12, 
    -4.61936e-13, -1.63522e-13, -2.538997e-13, -2.23481e-13, 1.057132e-12, 
    4.171802e-13, 1.650927e-12, 2.501693e-13, -4.810735e-13, -1.144154e-12, 
    6.094542e-13, -2.038689e-12, -3.831935e-13, 5.376064e-13, 2.755816e-12, 
    3.107237e-14, -1.739581e-13, 9.645063e-15, 3.483741e-13, 4.633793e-14, 
    -1.903339e-13, -8.75619e-13, -1.176961e-12, -3.738815e-13, -2.926132e-13, 
    8.788109e-13, 1.464021e-12, 1.345509e-11, -9.452794e-12, -1.19388e-12, 
    -4.912598e-13,
  5.629941e-13, 5.048462e-13, 5.445644e-13, 5.191403e-13, 1.356137e-13, 
    4.692358e-13, -4.859724e-13, 4.202194e-14, -7.106815e-13, -1.283224e-12, 
    -6.919465e-14, 6.632195e-13, -3.813339e-13, 7.385481e-13, -1.89268e-12, 
    7.171236e-13, 9.013151e-13, 5.838802e-13, 7.910929e-13, 1.424527e-12, 
    1.611683e-12, -1.736999e-12, -2.272571e-12, -1.619233e-12, -7.205625e-13, 
    -1.312006e-12, 2.669032e-12, 9.876544e-13, -1.67813e-12, 1.806388e-12, 
    -3.025885e-12, -5.273143e-12, -2.995659e-13, -7.436274e-13, 
    -2.151335e-12, -5.243306e-13, -7.181339e-13, -6.11608e-13, -1.165734e-14, 
    1.662032e-13, 4.194978e-13, 6.314393e-13, 8.117534e-13, 7.309531e-13, 
    -5.19873e-12, -2.08028e-13, -3.909373e-13, -2.061129e-12, -6.499634e-13, 
    1.482837e-11, 8.693532e-13, -3.032019e-13, -9.164558e-13, -2.288664e-12, 
    4.2569e-13, -2.986361e-13, -3.793632e-13, -3.175682e-13, -3.328726e-13, 
    -2.92464e-13, -1.901951e-12, -3.746087e-12, -4.401229e-12, 4.686917e-13, 
    5.722312e-13, -1.269596e-12, -1.300543e-12, 1.004447e-12, 3.546302e-12, 
    1.822903e-12, 7.405188e-14, -9.036938e-13, 1.805223e-13, -1.820488e-13, 
    9.366562e-13, -4.624634e-13, -6.456086e-13, -2.200393e-13, -9.28075e-13, 
    3.339273e-13, 1.317182e-12, -9.361262e-15, -4.575645e-13, 1.400852e-12, 
    -3.573253e-13, -5.298373e-12, -6.615097e-12, -5.385414e-13, 
    -3.324086e-13, -9.672541e-13, -1.252554e-12, 1.546485e-13, 3.040623e-14, 
    -2.250797e-12, 2.102984e-12, -8.787701e-12, 3.177292e-13, 1.64091e-13, 
    1.759612e-11, -3.946954e-13, -3.116035e-12, -2.627508e-12, 7.442276e-13, 
    2.075342e-12, 3.395617e-13, -3.415046e-13, -2.694234e-13, -9.759415e-13, 
    -9.842405e-13, -1.385309e-12, -8.271439e-13, -1.167871e-12, 1.132427e-14, 
    -8.363588e-13, 4.409556e-12, 2.900125e-12, 6.82147e-12, -2.897414e-12, 
    -1.97984e-13, -3.655132e-12,
  1.664224e-13, -3.614886e-13, 2.904899e-13, 3.625433e-13, -6.699086e-13, 
    1.772082e-12, -1.188938e-12, -2.274569e-12, -3.244904e-12, 2.838785e-12, 
    4.231837e-12, 8.521905e-12, 4.805267e-12, 6.106615e-12, -1.287193e-12, 
    2.407907e-13, 7.36966e-13, 8.670842e-13, -1.931164e-13, 1.412204e-12, 
    5.143108e-13, -3.885225e-13, -2.202682e-13, 9.056644e-13, -9.618972e-13, 
    -5.370038e-12, 2.834288e-12, 6.22008e-12, 1.806721e-12, -8.815171e-14, 
    -1.230072e-12, -2.087053e-12, -2.053968e-12, 3.576028e-13, -5.959067e-12, 
    -9.026557e-12, -1.403988e-13, -3.671854e-13, -3.960166e-12, 
    -5.260847e-13, -1.296108e-12, -5.816791e-12, 3.097897e-12, 6.710014e-13, 
    -3.235634e-12, 8.296419e-12, -3.849421e-13, 8.062995e-14, 1.299338e-12, 
    5.763903e-12, 1.700459e-12, -3.699263e-13, -3.858081e-13, 8.397705e-12, 
    -1.682279e-13, -4.27075e-13, -3.189671e-13, 8.521517e-14, -5.243861e-13, 
    5.696166e-12, -1.202322e-11, -6.226075e-12, -1.141687e-11, -4.55902e-13, 
    1.059342e-12, -1.531719e-11, -5.503098e-12, -4.76047e-12, -5.476841e-12, 
    -2.269851e-13, 2.414957e-12, -7.201517e-12, 3.943679e-12, -5.15088e-13, 
    -3.082562e-12, -5.991319e-13, -4.274775e-13, -1.800712e-12, 
    -8.514777e-12, -9.264589e-12, 3.046563e-12, -8.301425e-12, 1.423001e-12, 
    3.458955e-12, -9.801049e-13, -6.749046e-12, -1.657546e-11, -5.364598e-13, 
    -6.491535e-13, -8.820999e-13, -2.656153e-12, 5.6537e-13, -1.650208e-13, 
    -2.284612e-12, 5.440648e-13, -8.184564e-14, 1.082545e-12, 3.982925e-13, 
    1.360523e-11, 5.069589e-12, -4.050649e-12, -3.600158e-12, 7.753971e-13, 
    -8.052239e-14, 1.543932e-12, 4.652945e-13, -6.224465e-13, -1.222022e-12, 
    -4.250489e-13, -1.65773e-12, -8.26228e-13, -2.871037e-13, -3.470002e-13, 
    -4.765632e-13, -2.343237e-12, 6.145862e-12, 2.330351e-12, -1.473113e-12, 
    -1.142836e-14, -6.75926e-12,
  -2.341516e-12, -2.628009e-12, 1.564748e-12, -4.638345e-12, -3.393952e-12, 
    -4.198919e-12, -3.336498e-12, -4.757139e-12, 2.979311e-11, 3.049405e-11, 
    1.121864e-11, 5.444534e-13, -9.103607e-12, -4.595546e-12, 1.864664e-11, 
    1.639994e-12, -1.169442e-12, 2.248063e-12, 4.131251e-12, 1.471545e-12, 
    -1.594225e-12, -2.067402e-12, -2.630951e-12, 8.448797e-13, 1.221412e-12, 
    1.426825e-11, 1.482087e-11, 1.216965e-11, 1.907158e-11, 9.455214e-13, 
    -1.161049e-11, 8.311962e-12, -4.718448e-13, 6.096901e-12, -8.30408e-12, 
    -8.067935e-12, -2.133149e-12, -5.433987e-13, -1.786873e-10, 
    -2.611078e-13, 1.144096e-12, -9.640344e-12, 8.067297e-13, 2.178515e-12, 
    5.889456e-12, 3.529954e-13, -9.341139e-13, 3.565065e-13, -2.115008e-12, 
    -2.78132e-12, -1.608297e-13, -1.962985e-12, 1.876166e-12, 1.344166e-11, 
    -8.132439e-13, 1.601497e-14, -2.744416e-11, 3.121892e-13, -1.91534e-12, 
    8.525625e-12, -3.211564e-11, 1.766587e-12, -8.735124e-12, -1.85526e-12, 
    -2.423184e-12, 1.882344e-11, 2.470446e-11, -1.567851e-11, -2.174039e-12, 
    -1.171152e-11, -4.909406e-12, -2.462769e-11, 7.054357e-12, -2.434886e-12, 
    -6.288748e-13, -2.657874e-13, -2.764247e-13, 3.617939e-13, -1.620525e-11, 
    -1.52412e-11, -4.792361e-12, 5.534489e-13, 9.609258e-13, 1.55328e-11, 
    -1.67133e-12, -1.267431e-12, -4.804934e-12, 2.994327e-12, -5.732654e-13, 
    1.071643e-13, -9.544032e-13, -1.848538e-11, -3.394923e-13, -1.751499e-12, 
    1.837364e-12, -2.160794e-12, 7.807643e-13, 9.26581e-12, -2.061018e-12, 
    5.863932e-12, -1.249001e-14, -1.582887e-12, -1.507301e-13, -4.895761e-12, 
    -3.141931e-13, -1.016742e-12, -1.961764e-12, -3.102518e-13, 
    -9.947598e-13, -7.026046e-13, 4.20608e-13, -1.46716e-12, -5.812018e-14, 
    1.898315e-12, -2.727002e-11, 8.197782e-12, 2.78802e-12, -5.143452e-12, 
    4.307318e-14, 1.978973e-12,
  -1.174411e-11, -2.196254e-11, -2.122308e-11, -1.373202e-11, -8.002321e-12, 
    -1.085559e-11, 3.322342e-11, 3.348655e-11, 6.189049e-12, 6.599721e-12, 
    5.46696e-12, -2.789546e-12, -1.166844e-13, -5.494716e-12, 4.510003e-12, 
    1.519562e-12, -9.337103e-12, 2.791739e-12, 4.657177e-13, -9.376389e-13, 
    3.091472e-12, -1.908529e-12, 3.955614e-12, 2.034922e-11, 2.954875e-11, 
    4.649447e-11, 2.036693e-11, -1.968903e-11, 1.826245e-11, -3.446965e-12, 
    -4.693801e-12, -9.895529e-12, 1.738443e-12, -3.503697e-12, -7.865875e-12, 
    1.847483e-11, 2.396178e-12, -1.085139e-12, -1.290563e-10, 2.604417e-13, 
    -3.353984e-14, -7.225553e-12, 6.416243e-12, 5.767628e-12, 1.090317e-11, 
    -1.603662e-11, -6.713796e-13, -2.009712e-12, -6.596224e-12, 
    -5.174475e-12, -1.1732e-12, 9.321988e-13, 1.378175e-13, 1.039002e-12, 
    -5.429571e-12, 3.385625e-13, -2.424905e-11, 4.681089e-13, -1.278228e-12, 
    -8.452593e-12, -1.292244e-11, 2.211675e-12, -4.254486e-12, -7.165657e-12, 
    -1.093914e-12, -1.002032e-12, 1.599609e-12, 4.934664e-12, 2.340733e-11, 
    -9.241719e-12, 8.050782e-13, -9.731105e-13, 2.44299e-12, -1.730394e-12, 
    -3.589096e-12, -5.628831e-14, -3.963774e-13, -1.574435e-13, 
    -1.891811e-11, 3.804179e-13, -1.555506e-11, 1.66004e-11, -9.724999e-13, 
    3.912604e-11, -4.278744e-12, 4.924006e-12, -1.896039e-12, 6.224687e-12, 
    1.390893e-13, -1.042832e-12, -6.913914e-13, 3.61825e-12, -3.15234e-13, 
    3.826217e-13, -2.09871e-12, -1.989709e-12, -1.526346e-12, -3.677447e-12, 
    -1.07791e-11, 5.623224e-12, -4.708456e-12, -6.883626e-13, -4.390724e-13, 
    -1.035136e-11, -1.696088e-12, 4.686806e-13, 5.692891e-12, -1.180334e-12, 
    -3.561651e-12, -1.526224e-12, -6.826761e-13, 5.053291e-12, 5.853651e-12, 
    -2.83662e-12, -1.925299e-11, 1.732575e-12, 8.607559e-13, -3.998453e-12, 
    1.881134e-14, 8.956835e-12,
  -8.660295e-12, -5.765166e-12, -6.350476e-13, 1.696976e-12, 2.585293e-11, 
    4.210909e-12, 4.813649e-12, 1.015987e-11, 3.136658e-12, -3.554157e-12, 
    -8.895551e-12, 2.068457e-12, -1.132899e-11, -4.217737e-13, 5.505041e-13, 
    7.331358e-13, -6.944933e-12, 1.271844e-12, 4.405608e-12, 5.096645e-12, 
    5.674461e-12, -1.29563e-12, 5.310918e-12, 3.708317e-11, -8.874124e-12, 
    -2.753181e-11, -2.238981e-11, -1.586747e-11, -1.730849e-11, 6.647793e-12, 
    -1.540768e-12, -6.330431e-11, -3.610445e-13, -4.210521e-12, -5.96323e-12, 
    1.6321e-11, 1.389894e-12, -1.131907e-12, -2.82529e-11, -2.911837e-13, 
    -4.236844e-12, -3.667289e-12, 2.209205e-12, 1.428589e-12, 5.33823e-12, 
    9.833134e-12, -3.499701e-13, -3.977207e-12, 1.189677e-11, -2.913586e-12, 
    -1.230502e-12, -2.234052e-11, -1.052691e-12, 3.475997e-13, -4.885359e-12, 
    1.947331e-13, -2.110145e-12, 5.168588e-13, 3.964051e-14, -1.273889e-11, 
    1.965705e-12, -3.155254e-12, -6.708634e-12, -5.245881e-12, -4.401235e-12, 
    -3.439304e-12, 8.065937e-12, 1.154021e-12, 6.160517e-12, 3.237977e-11, 
    7.05902e-12, -6.935619e-12, -1.244183e-11, 9.546086e-12, -5.573442e-12, 
    8.354428e-14, -2.725112e-13, -5.385012e-11, -1.000278e-11, 9.743872e-13, 
    -1.545478e-11, 1.173666e-11, -3.662709e-12, -2.851869e-11, 4.215572e-12, 
    1.828343e-11, -7.573775e-12, 1.831507e-11, -7.511257e-13, -1.154687e-12, 
    -2.340517e-12, -1.442002e-12, 2.721712e-13, -6.311568e-12, -8.945844e-12, 
    -1.491401e-12, -1.199552e-12, -1.557848e-11, -1.235101e-11, 3.140954e-12, 
    -6.80983e-12, -5.032256e-12, -3.807163e-13, -1.253439e-11, 9.380829e-13, 
    1.662614e-12, 3.943512e-12, 2.363998e-12, -9.335588e-12, -3.764322e-12, 
    -7.87298e-12, 2.139566e-11, 9.6676e-12, 2.283029e-11, 3.63759e-12, 
    -1.10662e-12, 1.365574e-14, -3.487712e-12, 2.766731e-12, 3.85536e-12,
  5.557221e-12, 3.768746e-11, 5.167256e-11, 1.348843e-11, -5.625833e-11, 
    -4.732148e-11, -2.002781e-11, -2.511075e-11, -1.175188e-11, 
    -2.805789e-11, -1.731459e-11, 1.228811e-11, -5.715317e-12, -7.809864e-13, 
    -4.366285e-12, -2.663991e-12, -4.39685e-12, -8.780754e-13, 8.547052e-13, 
    1.049322e-11, 4.530487e-12, -9.627299e-13, 8.640588e-12, 1.094441e-11, 
    -5.032369e-11, -6.262135e-11, -1.151651e-11, 2.386891e-11, -7.07745e-12, 
    7.584011e-11, 5.153317e-11, 7.926254e-11, 4.895861e-12, 2.522482e-11, 
    -1.516642e-11, -2.488632e-11, -1.23318e-12, -6.651693e-13, 1.475131e-11, 
    -2.388273e-12, -1.282664e-11, -1.631284e-11, 5.888387e-12, -8.509339e-13, 
    -1.148048e-11, 4.618073e-11, 2.308709e-13, 1.301736e-14, 2.113423e-11, 
    4.256977e-13, 3.735671e-12, -7.85072e-12, -1.088246e-12, 1.165446e-12, 
    -4.712436e-12, 4.206635e-13, -1.469214e-12, 1.180184e-12, -1.384437e-12, 
    7.454773e-12, 7.548406e-12, -5.340173e-14, 1.759148e-13, -8.796919e-12, 
    -8.371803e-12, -3.91398e-12, 7.670498e-11, -8.598122e-12, 7.273959e-12, 
    1.101094e-10, 4.233669e-12, 1.701028e-11, -3.961886e-11, 4.436207e-11, 
    -3.993933e-12, 1.230127e-13, -1.929984e-13, -1.701128e-11, -2.605305e-13, 
    -2.667977e-12, -1.440534e-11, 3.601864e-12, -5.752898e-13, -6.423317e-11, 
    -1.164346e-12, 2.913247e-11, -5.436795e-11, 1.559053e-11, -1.427305e-12, 
    1.247696e-12, -5.088541e-12, 8.600898e-14, 2.412237e-12, -4.148387e-12, 
    -9.134693e-12, 7.389811e-13, -4.262002e-12, -3.034634e-11, -5.995204e-15, 
    -1.330158e-12, -5.487943e-12, -2.811005e-12, -8.806358e-13, 
    -6.124504e-12, 1.360084e-11, 3.137546e-12, -6.821044e-12, 3.282596e-12, 
    -1.758282e-11, -9.520162e-12, -1.465694e-11, 2.701506e-11, 4.528161e-11, 
    3.935885e-11, 1.671835e-11, -5.407119e-13, -1.954339e-13, -2.449192e-12, 
    5.674763e-12, -7.204515e-12,
  5.974699e-11, 7.565115e-11, 4.109457e-11, -3.219558e-11, -3.048128e-11, 
    -3.531475e-11, -2.893263e-11, -8.492684e-11, 3.743228e-12, -1.121356e-10, 
    -1.93443e-11, 2.969569e-11, -9.826362e-12, -5.286438e-12, -4.376355e-11, 
    -4.443856e-12, -3.627032e-12, -5.880796e-12, 1.235817e-11, 1.08159e-11, 
    1.250111e-12, -4.567902e-12, 4.180212e-12, 3.249623e-11, -1.50289e-10, 
    -6.227585e-11, -2.552747e-11, 3.732414e-11, 9.465206e-12, 5.180611e-11, 
    2.785661e-12, 5.790979e-11, 3.010825e-11, 1.794875e-11, -3.506384e-11, 
    5.77548e-11, -3.92697e-13, -2.309403e-13, 3.223932e-11, -2.303457e-12, 
    -8.469381e-12, -3.17133e-11, 5.82065e-12, -6.32449e-13, 3.030909e-13, 
    1.843925e-11, 1.983691e-12, 4.06164e-12, 5.777112e-12, 1.620371e-13, 
    2.086639e-11, 1.831268e-11, -8.458456e-13, 7.55418e-13, -1.998121e-12, 
    3.357314e-13, -1.093192e-10, 1.837874e-12, -1.751288e-12, 1.052768e-11, 
    1.39555e-12, -8.334777e-12, -1.792566e-12, -7.826739e-12, -9.165735e-12, 
    -4.340861e-12, 1.6493e-10, 2.779521e-11, -2.064326e-11, 9.164491e-11, 
    2.006539e-11, 3.082601e-11, 1.324385e-10, 5.087841e-11, 5.509815e-12, 
    6.794565e-14, 1.625089e-13, 1.086992e-11, 7.530837e-13, -6.306844e-12, 
    -1.380152e-11, -2.473799e-13, 1.736722e-12, -4.628153e-11, 3.392953e-12, 
    -8.932066e-11, -5.727829e-11, 8.937295e-12, -3.386683e-13, 4.260481e-13, 
    2.688405e-12, 7.176482e-13, 2.586376e-12, 8.954826e-12, -1.492506e-11, 
    3.570577e-12, -7.961076e-12, -2.119727e-11, 6.187939e-12, -1.450484e-12, 
    -5.092593e-12, 8.601252e-12, -1.064183e-12, 1.119105e-13, 2.505884e-11, 
    4.160472e-11, 1.215272e-11, -1.278422e-11, -2.208522e-11, -1.998324e-11, 
    -1.897671e-11, 8.227974e-12, 6.600076e-11, 4.51833e-11, 1.509914e-11, 
    2.237766e-13, -1.628558e-13, -1.141202e-12, 2.866075e-12, -9.3624e-12,
  1.440392e-10, 4.650502e-12, -1.403544e-11, -1.948997e-11, -2.908385e-11, 
    -3.493517e-11, -4.090572e-11, -1.252298e-10, -2.52794e-10, -1.513891e-10, 
    -4.25997e-11, 5.121348e-11, -9.424461e-12, -5.985434e-12, -5.743761e-11, 
    -6.108048e-12, -4.585288e-12, -1.736056e-12, 1.695172e-11, 1.015965e-11, 
    -5.235812e-13, -1.609624e-11, 2.926326e-11, 3.501222e-11, -2.415184e-10, 
    -9.500223e-11, -6.442402e-12, 3.367351e-11, 1.777467e-12, 1.525535e-11, 
    -4.536171e-11, 7.43805e-12, 1.04285e-10, -4.24405e-11, -7.248269e-11, 
    8.970247e-11, -1.159739e-13, -1.065814e-14, 1.117004e-10, 3.001821e-13, 
    -4.691847e-12, -2.289435e-11, 6.020184e-12, 2.173713e-13, 7.314438e-11, 
    -3.093348e-11, 8.109957e-12, 5.942469e-13, 3.611777e-13, -1.959127e-13, 
    2.241568e-11, -2.96474e-12, 4.790168e-13, 1.485034e-13, 1.046663e-13, 
    -1.117995e-13, -1.206701e-10, 1.610156e-12, 2.593126e-12, -5.134865e-12, 
    -4.763301e-12, -7.937029e-11, 1.903477e-11, -7.378498e-12, -6.772138e-12, 
    7.741274e-11, 6.804979e-11, 8.803025e-11, -1.433254e-11, 3.857004e-11, 
    7.786416e-11, 2.882847e-10, -1.14686e-11, 1.167728e-10, 2.813332e-11, 
    1.687539e-14, 2.589595e-13, 9.950263e-12, 6.470435e-13, -3.373346e-11, 
    -1.471334e-11, -2.116751e-12, -8.355538e-13, -3.727596e-11, 3.319323e-11, 
    -2.908527e-10, 1.010303e-10, 2.564837e-12, 3.746864e-13, -7.909229e-13, 
    2.193357e-12, 4.592326e-13, 1.20004e-12, -1.019633e-11, -2.639577e-11, 
    4.621214e-12, -9.132518e-12, -1.603229e-11, 1.30691e-11, 2.463807e-13, 
    1.500933e-11, 8.233969e-13, -6.942641e-13, 7.04159e-13, 3.153589e-11, 
    2.002865e-11, -2.185252e-11, -2.461809e-11, -2.370815e-11, -3.954947e-11, 
    -3.344858e-11, -1.703948e-11, 5.570744e-11, 3.709832e-11, 1.403389e-11, 
    1.670442e-13, 1.589284e-13, -2.273182e-14, 5.328793e-13, -1.884959e-11,
  4.644485e-11, -2.232636e-11, -2.064238e-11, -2.909295e-11, -7.489809e-11, 
    -6.137113e-11, -6.374479e-11, -1.746538e-10, -1.128038e-10, -2.47512e-10, 
    -1.833051e-10, 1.324711e-10, -8.841305e-11, 9.551693e-12, 6.094836e-11, 
    -8.375833e-12, -5.478507e-12, 1.293898e-11, 1.251182e-11, 1.176725e-11, 
    -9.15068e-12, -1.721712e-11, 5.441403e-11, 1.168288e-11, 5.855783e-11, 
    -2.674378e-10, 2.43896e-11, 6.647949e-11, 6.950596e-11, -2.701173e-12, 
    -1.273073e-10, -6.085576e-12, 2.149532e-10, -8.575207e-11, -2.808564e-10, 
    -5.028844e-11, -1.944178e-12, 8.126833e-14, 1.366918e-10, -8.169909e-13, 
    9.435341e-12, 1.11755e-12, 1.417644e-11, -4.926615e-16, 9.888068e-11, 
    -6.859779e-11, 2.058687e-11, 1.97975e-12, 8.794298e-13, -7.320533e-13, 
    -6.501799e-12, 2.817324e-11, 5.392531e-12, -2.302603e-13, -1.721956e-14, 
    -8.906209e-13, -1.762552e-10, 1.859002e-12, 1.856706e-11, -4.701495e-11, 
    -6.797007e-12, -1.773175e-10, 3.026046e-11, -5.207168e-12, 1.238565e-13, 
    6.456424e-10, -1.408096e-11, 1.47746e-10, -7.922329e-12, 5.223222e-11, 
    1.122153e-10, 5.435774e-10, -1.049394e-10, 1.89688e-10, 4.378031e-11, 
    1.401101e-13, 2.664535e-15, 5.511702e-12, -1.576006e-12, -1.200486e-10, 
    -1.498379e-11, -2.613087e-12, -4.962253e-12, -1.023959e-11, -3.25755e-11, 
    7.151548e-10, -1.543632e-11, 1.998179e-12, 1.5557e-14, -8.282264e-14, 
    1.502731e-11, 1.711031e-12, 4.08007e-13, -2.671237e-11, -4.314926e-11, 
    3.386713e-12, -1.379727e-11, 1.165668e-11, 1.537548e-11, 1.959455e-12, 
    3.572143e-11, 6.292775e-11, -4.374279e-14, 6.083745e-13, 2.259637e-11, 
    -9.731926e-11, -1.157778e-10, -7.262346e-11, -3.638356e-11, 
    -5.346812e-11, -4.275313e-11, -2.993628e-11, 1.886735e-11, -2.855272e-12, 
    1.828471e-11, -1.299849e-13, 7.944756e-13, 1.696004e-13, 1.184053e-13, 
    -1.558018e-10,
  3.159917e-12, -2.767764e-11, -5.391443e-11, -1.02091e-10, -1.051064e-10, 
    -1.083358e-10, -1.086413e-10, -1.934295e-10, -1.194709e-10, 
    -1.816887e-10, -1.124028e-10, 2.292244e-10, -2.276528e-10, 4.282508e-11, 
    2.733702e-11, -8.320766e-12, -4.086553e-12, 2.043987e-11, 2.522138e-11, 
    6.47904e-12, -2.2782e-11, -6.197043e-12, 5.381096e-11, 4.567702e-11, 
    4.093392e-12, -1.437137e-10, 5.337575e-11, 1.338571e-10, 1.269027e-10, 
    1.446376e-11, -2.752671e-10, -9.639511e-11, 2.385485e-10, -3.366447e-10, 
    -1.92488e-10, -1.236544e-11, -5.737855e-12, -3.974598e-14, 2.518943e-10, 
    -3.866285e-12, -1.635159e-11, 2.997491e-11, 1.579736e-11, -2.685782e-12, 
    1.893621e-10, -7.962719e-11, 3.781531e-11, 1.461031e-11, 1.070388e-12, 
    -1.937284e-12, -2.581491e-11, 4.577028e-11, 1.779461e-11, 1.876321e-12, 
    1.806333e-13, -5.833112e-13, 4.320933e-10, 3.364464e-12, 4.88289e-11, 
    -1.024013e-10, -3.496092e-12, -1.200056e-10, 6.230194e-11, 4.766099e-12, 
    1.765854e-11, 1.504661e-10, -2.195713e-10, 2.6231e-10, 2.901834e-11, 
    8.124235e-11, 7.906276e-11, 7.247596e-10, -2.458711e-10, 1.580325e-10, 
    4.980181e-11, -1.023626e-13, -9.769963e-15, 1.08924e-11, -7.723089e-12, 
    -7.108469e-11, -1.538258e-11, -5.198819e-12, -8.255396e-12, 
    -8.913981e-12, 5.759904e-11, 3.550775e-10, 4.765766e-11, 6.339596e-12, 
    -1.29291e-12, -4.891643e-13, 4.174217e-12, -1.28296e-11, 7.460699e-13, 
    -2.972009e-11, -8.395351e-11, -8.606005e-13, -2.718736e-11, 
    -9.604073e-11, 1.119971e-11, 5.467582e-12, 4.132139e-11, 4.668886e-10, 
    3.506639e-13, 4.573009e-13, -2.836176e-12, -1.2226e-11, -2.094442e-10, 
    -2.011993e-10, -4.615974e-11, -5.692535e-11, -4.28193e-11, -3.965739e-11, 
    -3.305201e-11, -6.241963e-11, 1.917555e-11, -1.292744e-13, 1.651901e-12, 
    -6.386558e-14, -4.611866e-13, -3.89295e-10,
  1.421419e-11, -3.838729e-11, -1.124933e-10, -1.581617e-10, -1.5001e-10, 
    -1.424871e-10, -1.71821e-10, -1.847458e-10, -2.810634e-10, 1.604146e-10, 
    1.338374e-11, 5.575724e-10, -2.398315e-10, 9.690893e-11, -3.485678e-11, 
    -3.615375e-12, -1.427347e-12, 1.129341e-11, 5.300238e-11, -1.935452e-11, 
    -2.902678e-11, 6.759704e-12, 3.467959e-11, -7.318612e-11, -6.39311e-10, 
    -7.635814e-10, 5.310663e-11, 2.126839e-10, 3.043217e-10, 5.310485e-11, 
    -5.18088e-10, -1.576359e-10, 2.883513e-10, -1.838907e-11, 1.82222e-10, 
    1.10745e-10, -9.835732e-12, -2.078338e-13, 5.350962e-10, -4.461098e-12, 
    -4.528879e-11, 2.615752e-11, 3.75322e-12, -7.394904e-12, 3.330658e-10, 
    -1.642004e-10, 5.109313e-11, 9.536594e-12, 1.083711e-12, -4.264533e-12, 
    2.542966e-12, 8.163226e-11, 4.955862e-11, 4.703748e-12, 3.411027e-12, 
    9.547918e-15, 1.349265e-10, 7.001555e-12, 7.943801e-11, -1.147389e-10, 
    -7.081669e-12, 7.680057e-11, 1.507112e-10, 1.34786e-11, 1.973564e-11, 
    1.822478e-10, 7.612022e-11, 2.73066e-10, 6.093415e-11, 1.502947e-10, 
    4.261902e-11, 1.614736e-09, 7.202039e-11, 1.3034e-10, 5.820433e-11, 
    -1.637135e-12, 2.271516e-13, 2.764944e-11, -1.000162e-11, 7.119527e-11, 
    -1.903255e-11, -4.051448e-12, -7.551959e-12, -1.033773e-11, 
    -2.868839e-11, 1.003196e-09, 3.203871e-10, 1.503397e-11, -6.396675e-12, 
    -1.608647e-11, 4.662026e-11, -1.512612e-12, -2.624567e-13, -1.550169e-11, 
    -8.209367e-11, -1.018576e-11, -4.955969e-11, -2.108627e-10, 8.607115e-12, 
    8.807488e-12, 1.88211e-10, 7.779928e-10, 1.692646e-12, 1.905698e-12, 
    2.350897e-11, 2.732177e-10, -1.739162e-10, -3.55554e-10, -5.087242e-11, 
    -4.394907e-11, -3.811551e-11, -3.318257e-11, -7.226775e-11, -1.18906e-10, 
    2.162515e-11, 2.722267e-14, 1.857736e-12, 2.953193e-13, -1.963263e-12, 
    -2.928948e-10,
  2.265743e-11, 6.597034e-11, -1.093525e-10, -3.381668e-10, -3.601084e-10, 
    -2.16124e-10, -2.602523e-10, -1.511058e-10, -5.653469e-10, 2.468532e-10, 
    8.482637e-11, -1.044741e-09, 1.513225e-10, 1.524398e-10, -3.772982e-11, 
    4.134293e-12, 3.067058e-12, -5.672796e-12, 7.505374e-11, -5.088019e-11, 
    -3.348077e-11, 4.24194e-12, 6.247447e-12, -3.101253e-10, -1.295136e-09, 
    -1.182908e-09, -1.640981e-10, 5.530136e-10, 5.752767e-10, -2.312106e-11, 
    -1.07484e-09, -4.674305e-10, 3.399041e-10, 5.439453e-10, 5.562946e-10, 
    4.670131e-10, -1.31628e-11, 1.554312e-14, 8.509957e-10, -1.800995e-11, 
    4.285816e-11, -5.989875e-12, -3.023803e-12, -1.160408e-11, 3.509193e-10, 
    -4.589076e-10, 6.083578e-11, -5.915535e-11, 1.843858e-13, -7.719714e-12, 
    4.587086e-11, 3.36227e-10, 1.266706e-10, -4.757084e-12, 9.699841e-12, 
    -3.28626e-14, -1.40842e-10, 1.80453e-11, 1.148264e-10, 5.170819e-11, 
    -7.885248e-12, 1.639435e-10, 1.216591e-10, 8.165557e-12, 6.603074e-12, 
    7.149836e-11, -1.833556e-11, 7.318288e-10, 1.623519e-10, 1.649543e-10, 
    5.126921e-11, 3.193435e-09, 2.720935e-10, 3.155129e-10, 9.636487e-11, 
    -4.186873e-12, 4.856116e-13, 4.648726e-11, -2.766232e-12, 2.404708e-10, 
    -3.402345e-11, -8.731682e-13, -2.133405e-12, -2.758682e-12, 4.777867e-11, 
    9.359233e-10, 3.758132e-10, 2.892619e-11, -2.707351e-11, -7.526069e-11, 
    1.736158e-10, 1.356135e-10, -4.440448e-12, 2.881429e-12, -6.865619e-11, 
    -2.268799e-11, -7.333192e-11, -3.096012e-10, 6.888712e-12, 1.073843e-11, 
    6.004939e-10, 6.595783e-10, 4.818923e-12, 5.708989e-12, 9.7236e-11, 
    4.170282e-10, -4.103917e-11, -3.99627e-10, -8.075318e-11, -2.664891e-11, 
    -3.045919e-11, -2.462741e-11, -1.306866e-10, -1.816769e-10, 1.783818e-11, 
    6.799894e-13, 7.929213e-13, 1.226963e-12, -4.518275e-12, 7.320367e-11,
  3.701928e-12, 1.867111e-10, 2.492637e-10, -5.828227e-11, -5.551328e-10, 
    -4.9228e-10, -3.46521e-10, -1.720579e-10, -4.866969e-10, 6.006111e-10, 
    -6.672618e-10, -8.977405e-10, 3.591101e-10, 2.037126e-10, 4.805223e-11, 
    1.574989e-11, 1.675584e-11, -2.715517e-11, 8.05076e-11, -6.98428e-11, 
    -4.155432e-11, -1.001688e-11, 4.583001e-13, -4.459224e-10, -1.430575e-09, 
    -1.731228e-09, -2.909637e-10, -9.44862e-11, 5.620198e-10, -2.57101e-10, 
    -1.67198e-09, 5.259384e-10, 6.867857e-10, -8.286811e-10, 3.786234e-10, 
    6.471712e-10, -1.853859e-11, 1.745493e-12, 1.111538e-09, -9.499228e-11, 
    -5.773764e-11, -6.659029e-11, 1.62137e-12, -1.356515e-11, 6.406271e-10, 
    -8.211849e-10, 8.242029e-11, -1.237526e-10, 3.850431e-12, -1.389056e-11, 
    4.652789e-11, 8.539303e-10, 2.822629e-10, -3.22359e-11, 8.902257e-12, 
    3.481659e-13, -8.918786e-10, 3.5479e-11, 2.161965e-10, 2.685379e-10, 
    1.793943e-11, 1.349694e-10, 1.2807e-10, -3.690204e-12, -4.966339e-12, 
    -2.273843e-10, -6.7649e-10, 4.969429e-10, 3.778524e-10, 2.289688e-10, 
    1.544755e-10, 5.165251e-09, 2.34941e-10, 7.365255e-10, 1.501434e-10, 
    -5.433876e-12, 5.482281e-13, 4.523137e-11, 6.157475e-12, 4.359766e-10, 
    -7.134915e-11, -3.675233e-11, 6.735057e-12, 1.923084e-11, 8.029133e-12, 
    -6.804584e-10, 8.14353e-11, 3.675105e-11, -8.899437e-11, -1.657394e-10, 
    5.514362e-10, 4.420311e-10, -7.264855e-12, 6.10374e-11, -2.835083e-10, 
    -2.732303e-11, -8.967049e-11, -2.876757e-10, 2.181366e-12, 1.257163e-11, 
    1.178812e-09, 4.517039e-10, 8.406054e-12, 6.46494e-12, 1.371312e-10, 
    4.896474e-10, 2.217533e-10, -7.283987e-10, -5.61327e-10, -6.247625e-11, 
    -2.019718e-11, -4.23217e-11, -1.987672e-10, -3.024727e-10, -4.583001e-13, 
    2.241229e-12, -2.1525e-12, 2.227774e-12, -5.819456e-12, 2.857714e-10,
  4.423129e-12, -3.538503e-12, 3.487699e-11, 6.028209e-10, 3.699476e-10, 
    -1.76307e-10, -4.542713e-10, -3.288569e-10, -1.788045e-10, 4.057767e-10, 
    -1.075176e-09, 6.044942e-11, 4.739e-10, 2.870628e-10, 2.48999e-10, 
    1.938289e-11, 4.045973e-11, -4.15632e-11, 7.562617e-11, -7.516476e-11, 
    -5.069722e-11, -1.072209e-11, 4.330758e-11, -2.735305e-10, -1.702031e-09, 
    -2.518259e-09, -3.862226e-10, -6.296581e-10, -5.483045e-10, 
    -5.728644e-10, -2.541057e-09, 6.526264e-10, 1.648083e-09, -1.223583e-09, 
    1.9919e-10, -5.917755e-11, -2.846825e-11, 5.373479e-12, 1.795016e-09, 
    -2.422667e-10, -3.130573e-10, -1.89992e-10, 3.182343e-12, -1.599415e-11, 
    6.02089e-10, -9.681642e-10, 1.305214e-10, -1.550671e-11, 1.87832e-11, 
    -2.785994e-11, -9.065948e-11, 8.817764e-10, 5.121425e-10, -5.822827e-11, 
    -8.293632e-12, 1.538325e-12, 5.34893e-10, 4.470557e-11, 5.231279e-10, 
    -2.330118e-10, 5.091749e-11, 5.419309e-11, 2.154366e-11, -5.410073e-12, 
    -8.517987e-12, -8.943779e-10, -9.029719e-10, -4.22574e-10, -2.7703e-10, 
    4.48118e-10, 3.987317e-10, 5.664099e-09, -7.876011e-10, 1.065366e-09, 
    2.351456e-10, -3.385736e-12, 9.237056e-14, 2.92788e-11, 1.296359e-11, 
    5.571508e-10, -1.361595e-10, -1.039666e-10, 9.922729e-12, -5.232614e-10, 
    -1.674607e-10, -3.568392e-09, -3.019451e-11, 5.704948e-11, -1.852365e-10, 
    -3.262901e-10, 1.156568e-09, 8.131117e-10, -2.375877e-12, 1.069342e-10, 
    -9.074341e-10, -2.145377e-11, -9.389467e-11, -5.605116e-11, 
    -1.598721e-13, 1.387406e-11, 1.696257e-09, 3.35701e-10, 9.793277e-12, 
    -7.41962e-12, 1.126459e-10, 4.992451e-10, 9.240892e-10, -1.375216e-09, 
    -1.957147e-09, -4.576073e-10, 8.778756e-12, -7.229062e-11, -3.702318e-10, 
    -5.928271e-10, -3.350564e-11, 6.771472e-12, -1.847411e-13, 3.359091e-12, 
    -5.197398e-12, 3.033804e-10,
  7.460343e-11, 2.518696e-10, -4.591527e-11, 3.06013e-10, 6.220873e-10, 
    7.440484e-10, -2.463452e-10, -4.83162e-10, -4.304965e-10, 3.764455e-10, 
    -2.173195e-10, 6.83869e-10, 5.992469e-10, 4.714309e-10, 4.819967e-10, 
    -3.034053e-11, 6.249365e-11, -2.215295e-11, 6.867795e-11, -7.2788e-11, 
    -6.108891e-11, -9.162449e-12, 4.14353e-11, -8.33289e-11, -1.319176e-09, 
    -3.090996e-09, -7.334542e-10, 7.560885e-11, -2.322334e-09, -9.629559e-10, 
    -3.843205e-09, 3.117755e-10, 1.933618e-09, -1.993286e-09, 1.876295e-10, 
    -1.645859e-09, -3.916476e-11, 9.758416e-12, 1.649784e-09, -3.927248e-10, 
    -4.844957e-10, -3.221352e-10, -1.815614e-11, -2.501321e-11, 
    -1.685393e-09, -8.914327e-10, 2.521787e-10, 8.969447e-11, 2.679101e-11, 
    -3.444423e-11, -1.472729e-10, 5.100631e-10, 7.626216e-10, -1.088765e-10, 
    -8.981082e-12, 2.184919e-12, 3.643315e-09, 3.954206e-11, 1.067472e-09, 
    2.6643e-10, 9.080381e-11, -3.79039e-11, 5.79103e-10, 1.506635e-11, 
    5.901768e-12, -1.286928e-09, -1.176165e-09, -1.984777e-09, -7.708714e-10, 
    1.311523e-09, 1.168697e-09, 3.044068e-09, -4.782059e-10, 8.143495e-10, 
    3.221562e-10, 4.721556e-12, -1.167066e-12, 5.629008e-11, 3.799974e-11, 
    6.571632e-10, -2.083187e-10, -2.569513e-10, -4.002132e-12, -1.172566e-09, 
    -7.738521e-11, -1.452548e-09, -8.190071e-11, 1.075335e-10, -2.591135e-10, 
    -4.54401e-10, 1.306798e-09, 9.710192e-10, 1.55973e-11, 6.393357e-11, 
    -2.34855e-09, 6.326673e-12, -1.286288e-10, 4.875531e-10, -1.964651e-12, 
    1.352092e-11, 1.692626e-09, 2.996963e-10, 9.03988e-12, -2.835909e-11, 
    -3.936407e-12, 3.588099e-10, 1.013902e-09, -9.074874e-10, 3.907132e-10, 
    -6.839009e-10, -6.495071e-11, -6.550138e-11, -6.848992e-10, 
    -1.065715e-09, -5.883649e-11, 1.245084e-11, 1.78515e-11, 3.875122e-12, 
    -3.227196e-12, 1.549374e-10,
  1.86553e-10, -9.103331e-10, -6.370513e-10, 3.965255e-10, 3.525571e-10, 
    7.696741e-10, 4.098766e-10, -4.556426e-10, -1.356163e-09, 3.302958e-10, 
    6.681304e-10, -1.28999e-10, 6.685426e-10, 7.065069e-10, 9.332339e-10, 
    -1.486185e-10, 5.092815e-11, 1.535838e-11, 9.539036e-11, -6.790657e-11, 
    -7.911183e-11, 8.39151e-12, -1.104823e-10, -1.77333e-09, -8.745502e-10, 
    -2.660904e-09, -1.803343e-09, 1.952628e-09, -8.401955e-10, -2.996309e-09, 
    -5.422677e-09, -1.390461e-10, 4.617036e-10, -3.54062e-09, 1.903615e-10, 
    -2.058123e-09, 3.15552e-11, 1.209433e-11, -2.569109e-09, -5.409909e-10, 
    -7.582912e-10, -3.058958e-10, -3.796785e-11, -4.314071e-11, 
    -3.083358e-09, -6.942074e-10, 5.406982e-10, -2.427907e-10, 1.905533e-11, 
    -4.377476e-11, 1.259473e-10, -4.827427e-11, 7.307946e-10, -1.397467e-10, 
    5.793978e-11, -2.096101e-13, 5.892332e-09, 4.967973e-11, 1.638033e-09, 
    8.620962e-10, 1.478355e-10, -1.025242e-10, 4.989289e-10, 3.64011e-11, 
    4.322658e-11, -2.739661e-09, -3.874149e-09, -6.185253e-09, -2.785683e-10, 
    1.560721e-09, 2.347626e-09, -2.914078e-10, -2.957634e-10, 3.487344e-11, 
    6.335085e-10, 2.756195e-11, -4.928502e-12, 1.131326e-10, 9.242562e-11, 
    9.979431e-10, -2.492051e-10, -5.291276e-10, 6.309619e-12, -1.113634e-10, 
    -2.506653e-10, 1.457245e-09, 6.688623e-10, 1.663878e-10, -3.180165e-10, 
    -6.20755e-10, 1.131468e-09, 7.172901e-10, 5.215206e-11, 3.677343e-11, 
    -2.79227e-09, 4.345111e-11, -2.706983e-10, 1.364342e-09, -4.973799e-12, 
    1.693507e-11, 1.096005e-09, 2.57653e-10, 7.521095e-12, -4.352074e-11, 
    -2.481428e-10, 3.126388e-12, 5.325802e-10, -1.438409e-09, 1.983693e-10, 
    -8.675087e-10, 3.645084e-11, -4.758505e-11, -8.780887e-10, -1.29117e-09, 
    -1.948308e-11, 2.154792e-11, 8.301981e-11, 1.334488e-13, -3.759215e-12, 
    5.318412e-11,
  2.364935e-10, -4.026621e-09, -7.940148e-09, -1.4923e-09, 5.764882e-10, 
    1.18245e-10, 1.448225e-09, -5.538325e-11, -2.572182e-09, 1.277666e-09, 
    1.940176e-09, -1.835918e-09, 1.428941e-09, 8.724292e-10, 2.148948e-09, 
    -5.018087e-10, -1.482995e-10, 7.968737e-12, 2.197744e-10, -5.056577e-11, 
    -1.060023e-10, -7.336354e-12, -3.210125e-10, -3.039322e-09, 
    -7.713261e-10, -8.522854e-10, -3.818986e-09, 2.691419e-09, 3.086136e-10, 
    -6.502052e-09, -6.446275e-09, 2.190141e-10, -2.393143e-10, -4.363816e-09, 
    1.925677e-10, -3.221079e-09, 2.557137e-10, 1.224798e-11, -1.313058e-09, 
    -7.742308e-10, -1.061634e-09, -9.064038e-11, 4.034106e-11, -9.818568e-11, 
    -5.409678e-09, -2.485798e-10, 1.05619e-09, 1.481588e-10, 1.795897e-11, 
    -2.081091e-11, -1.05782e-10, 4.397904e-11, -1.729866e-10, -5.786447e-11, 
    7.759163e-11, -8.004264e-12, 3.901132e-09, 1.090562e-10, 2.070637e-09, 
    1.630715e-09, 1.642597e-10, -2.996252e-10, 1.065068e-10, -7.356249e-12, 
    5.852527e-11, -7.417842e-09, -1.209323e-08, -1.100505e-08, 3.744898e-09, 
    -5.852065e-10, 6.010588e-10, -2.004246e-09, 1.488409e-10, -3.86553e-10, 
    9.192412e-10, 5.67546e-11, -1.137757e-11, 1.406804e-10, 8.913688e-11, 
    1.457732e-09, -2.437197e-10, -1.057496e-09, 8.478551e-11, 7.968701e-10, 
    -3.794618e-10, 1.412356e-09, 9.441941e-10, 1.983089e-10, -4.432381e-10, 
    -5.530474e-10, 1.013714e-09, 2.721798e-10, 9.410073e-11, 9.299228e-11, 
    -1.97193e-09, 9.990871e-11, -4.817799e-10, 2.121748e-09, -1.464073e-11, 
    1.130829e-11, 5.834622e-11, 1.566569e-10, 5.35838e-12, -5.409095e-11, 
    -4.976677e-10, -5.608065e-10, -9.911005e-11, -3.538137e-09, 2.700169e-10, 
    -1.922107e-09, 2.639347e-10, -2.433787e-10, -9.084182e-10, -1.361474e-09, 
    1.05711e-10, 3.078284e-11, 1.766818e-10, -1.381073e-11, -1.770939e-11, 
    -1.199716e-10,
  1.830536e-10, -8.600054e-11, -7.52102e-09, -7.133149e-09, -3.403013e-09, 
    7.218439e-10, 1.479709e-09, 7.90795e-10, -2.072323e-09, 3.03017e-09, 
    5.538613e-09, -5.440992e-09, 1.172044e-09, 9.805099e-10, 2.606004e-09, 
    -8.954494e-10, -4.24496e-10, -7.701928e-11, 3.575202e-10, -2.837552e-11, 
    -9.572076e-11, -6.360423e-11, -3.046914e-10, -1.887098e-09, 4.099622e-09, 
    6.758718e-10, -3.536652e-09, 4.493319e-09, 1.463111e-09, -8.229971e-09, 
    -6.680917e-09, 5.723457e-10, -4.350191e-10, -3.22208e-09, 8.242651e-11, 
    -4.446232e-09, 4.146706e-10, 2.74909e-11, -1.270418e-09, -7.012609e-10, 
    -1.121224e-09, 9.208989e-11, 2.024372e-10, -3.888938e-10, -5.312256e-09, 
    5.199787e-10, 1.831939e-09, 3.671339e-10, 9.363319e-11, -9.003465e-12, 
    -2.576517e-10, -2.159695e-11, -3.128875e-11, -2.025921e-10, 
    -9.840697e-11, -1.715605e-11, 7.095014e-09, 2.12777e-10, 2.199977e-09, 
    9.78325e-10, 1.308429e-10, -6.120437e-10, -2.781775e-12, -5.277421e-10, 
    3.01533e-11, -1.170951e-08, -9.832529e-09, 2.196575e-09, -6.908039e-10, 
    8.609113e-10, -2.294765e-09, 8.172272e-10, 4.415348e-10, 7.387122e-10, 
    5.472508e-10, 4.786571e-11, -8.306245e-12, 1.590159e-10, -7.529231e-11, 
    7.754046e-10, -4.051337e-10, -1.851245e-09, 2.617604e-10, 2.051966e-09, 
    4.939018e-10, 5.431282e-10, 1.307175e-09, 1.903011e-10, -7.392116e-10, 
    -1.259544e-10, 1.112912e-09, -1.747956e-10, 1.201563e-10, 7.591225e-11, 
    -1.646409e-09, 2.048573e-10, -5.573263e-10, 2.330101e-09, -3.583622e-11, 
    -3.630874e-13, -9.622845e-10, -7.270362e-11, 1.27276e-12, -2.154454e-11, 
    -6.581438e-10, -1.888363e-09, -2.10245e-09, -3.081649e-09, -3.830785e-10, 
    8.854677e-10, 1.439577e-09, -4.766001e-10, -1.137021e-09, -1.344713e-09, 
    3.099423e-10, 2.954934e-11, 1.428937e-10, -3.750156e-11, -5.601031e-11, 
    -4.333565e-10,
  -1.710596e-10, 3.08837e-09, -1.222368e-08, -1.391346e-09, -1.017505e-08, 
    -1.14456e-09, 1.757137e-10, 2.235634e-09, 1.284871e-09, 4.207617e-09, 
    7.281681e-09, -1.618208e-09, 1.620361e-09, 6.237251e-10, 2.155911e-09, 
    -6.005487e-10, -4.663129e-10, -3.197762e-10, 6.582432e-10, -1.429221e-10, 
    -1.310134e-10, -1.593499e-10, -2.29921e-10, -7.233787e-10, 1.305933e-08, 
    3.887504e-09, -3.091618e-09, 9.022056e-09, 3.640491e-09, -9.38822e-09, 
    -4.882867e-09, -6.59572e-10, 2.813788e-09, -3.31308e-09, 5.935519e-11, 
    -3.763962e-09, 5.114906e-10, 4.664713e-11, 2.945693e-09, -9.821466e-11, 
    -7.191325e-10, -2.071836e-10, 9.725802e-10, -6.928587e-10, -7.158754e-10, 
    1.040586e-09, 2.849017e-09, 4.826539e-10, -3.398789e-10, 1.911893e-11, 
    -4.009877e-10, -5.330101e-10, 6.927614e-10, 2.58165e-10, -2.396661e-10, 
    -2.119194e-11, 1.43235e-08, 3.294069e-10, 1.3488e-09, 8.450023e-10, 
    9.482548e-11, -6.886758e-10, 2.911449e-11, -3.724086e-09, 1.975238e-11, 
    -1.45934e-08, -6.089142e-09, 1.702784e-09, -3.246626e-09, 4.023786e-09, 
    -1.68659e-09, 5.335192e-09, 8.536283e-10, 7.241105e-10, 3.488772e-13, 
    3.687362e-11, 8.14282e-12, -5.272582e-11, 8.573408e-12, 4.937917e-11, 
    -1.408626e-09, -2.340643e-09, 6.161223e-10, 7.158103e-09, 6.602754e-10, 
    4.643397e-12, 8.988188e-10, 1.629523e-10, -1.313362e-09, -7.493739e-11, 
    8.003092e-10, 2.196821e-10, 1.204619e-10, 9.978507e-11, 8.838121e-10, 
    2.979441e-10, -4.381725e-10, 1.929077e-09, -8.50271e-11, -1.961738e-11, 
    -2.603038e-10, -6.394973e-10, -1.423928e-11, 6.314593e-11, -1.184805e-09, 
    -3.535821e-09, -5.461221e-09, -6.244523e-09, -5.282391e-09, 4.93905e-09, 
    4.711449e-09, -8.708305e-10, -1.484739e-09, -1.35886e-09, 4.652456e-10, 
    3.887379e-12, -1.888125e-10, -4.146727e-11, -8.223111e-11, -6.232774e-10,
  -9.445174e-10, 2.966651e-09, -4.641215e-09, -1.056006e-08, -4.946294e-09, 
    -8.461974e-09, -5.50564e-10, 2.603876e-09, 2.997062e-09, 4.344535e-09, 
    7.30963e-09, 5.317808e-09, 1.503246e-09, -3.498499e-10, 1.02613e-09, 
    -5.442402e-10, -2.728555e-10, -3.021299e-10, 1.259796e-09, -4.295231e-11, 
    -2.065761e-10, -2.949108e-10, -1.189804e-10, 4.659384e-10, 1.510062e-08, 
    7.184944e-09, -2.999521e-09, 1.31763e-08, 3.378737e-09, -1.128692e-08, 
    -2.458542e-09, 5.151648e-10, 6.595052e-09, -5.003393e-09, -1.066169e-10, 
    -3.64907e-09, 3.594934e-10, 1.611866e-11, 7.409874e-09, 1.650378e-10, 
    5.565965e-11, -8.621512e-10, 3.413824e-09, -9.554393e-10, 3.27784e-09, 
    1.720103e-09, 3.571692e-09, 5.344205e-10, -5.221935e-10, -1.393232e-10, 
    -5.215277e-10, -1.485326e-09, 2.065492e-09, 1.084217e-10, -1.034259e-10, 
    -3.060308e-11, 1.98749e-08, 4.435478e-10, 7.782873e-10, 2.416556e-11, 
    1.48809e-10, -6.830376e-10, -2.484697e-10, -9.029903e-09, -5.492495e-12, 
    -1.415442e-08, -4.658894e-09, -1.221316e-09, 1.200274e-08, 5.336595e-09, 
    -1.06116e-09, 1.312741e-08, 1.730676e-09, -5.558221e-10, 8.715514e-12, 
    6.740919e-11, 7.140954e-12, -8.15966e-10, 1.854076e-10, -2.291991e-09, 
    -2.038085e-09, -3.01374e-09, 1.163748e-09, 8.491689e-09, 2.035272e-09, 
    -9.122303e-10, 6.776233e-10, 8.127898e-11, -2.001833e-09, -8.704859e-11, 
    -1.463214e-09, 2.073038e-09, 8.488144e-11, 2.350092e-10, 3.19644e-09, 
    4.257757e-10, -3.270387e-10, 2.343022e-09, -2.00977e-10, -2.774669e-11, 
    4.002843e-10, -1.363295e-09, -3.281286e-11, 2.165699e-10, -2.179554e-09, 
    -2.48918e-09, -4.729777e-09, -8.492329e-09, -5.152579e-09, 3.710674e-09, 
    9.966008e-09, -9.604335e-10, -1.805752e-09, -1.62499e-09, 2.799467e-10, 
    -1.425491e-11, -7.343175e-10, 8.321344e-12, -9.911716e-11, -6.97618e-10,
  -2.069527e-09, 1.303704e-09, 1.864464e-10, -7.797951e-09, -3.228621e-09, 
    -9.652183e-09, -8.469669e-11, 2.239176e-09, 3.12744e-09, 4.616624e-09, 
    5.327905e-09, 1.173632e-08, 1.251806e-09, -2.235765e-09, 1.432909e-09, 
    -6.605374e-10, -6.315133e-10, -2.58126e-10, 1.520942e-09, 2.50111e-10, 
    -3.228706e-11, -5.478284e-10, -6.804157e-11, 1.273975e-09, 7.224855e-09, 
    5.966228e-09, -1.280398e-10, 1.222634e-08, 5.254009e-09, -1.385001e-08, 
    -1.38499e-09, 3.097256e-09, -1.650392e-09, -4.087696e-09, 1.089688e-10, 
    -3.625757e-09, 4.223182e-11, -8.504486e-11, 1.315146e-08, -7.969714e-11, 
    6.697632e-10, -1.127574e-09, 7.739693e-09, -1.368997e-09, 5.380002e-09, 
    2.20399e-09, 3.750685e-09, 6.58531e-10, -9.331473e-10, -2.984368e-10, 
    -5.433485e-10, -7.248104e-10, 4.164065e-09, -1.839737e-10, -3.337796e-10, 
    -7.078427e-11, 2.598637e-08, 5.537004e-10, 4.40042e-10, -2.129184e-09, 
    1.303988e-10, -1.522096e-09, -9.960388e-10, -1.310481e-08, -9.784913e-10, 
    -9.724204e-09, -4.6455e-09, -9.921166e-10, 1.93894e-08, 5.533764e-09, 
    -1.591445e-09, 2.333766e-08, 1.42694e-09, -1.662499e-09, -2.782556e-09, 
    1.701608e-10, -5.396572e-12, -2.044281e-09, 3.77441e-10, -1.372229e-09, 
    -1.107921e-09, -4.876727e-09, 1.76972e-09, 2.491845e-09, 2.006232e-09, 
    -7.734968e-10, 1.637147e-09, -5.192646e-11, -2.415193e-09, -7.847802e-10, 
    -4.925653e-09, 6.037573e-09, -3.183231e-12, -2.506101e-09, 3.310873e-09, 
    6.311097e-10, -3.851483e-10, 3.834828e-09, -2.929994e-10, -3.175273e-11, 
    2.020982e-09, -9.926087e-10, -2.971312e-11, 3.228582e-10, -2.105821e-09, 
    -6.109815e-10, -3.429335e-09, -5.826479e-09, -2.895888e-09, 9.522267e-09, 
    1.502161e-08, -1.544038e-09, -2.674284e-09, -2.255462e-09, -3.019522e-10, 
    -4.287415e-11, -2.770975e-10, 5.888356e-11, -9.159784e-11, -7.401297e-10,
  -2.981295e-09, 1.96053e-09, 1.067184e-08, 1.843944e-09, -1.740858e-09, 
    -2.586006e-09, -2.353175e-09, 2.046789e-09, 3.264091e-09, 3.780229e-09, 
    4.363301e-09, 1.651838e-08, 1.604946e-09, 2.029026e-10, 1.325589e-10, 
    -3.134346e-10, -1.352973e-09, -1.058439e-09, 1.188322e-09, 3.197727e-09, 
    -8.135714e-10, -9.424923e-10, -7.997869e-11, -2.448814e-10, 
    -5.481127e-10, 1.245022e-08, 1.458346e-09, 5.35448e-09, 1.656232e-08, 
    -2.26774e-08, -6.336336e-09, 5.005347e-09, 2.008932e-09, -4.420315e-09, 
    -2.131344e-10, -1.688278e-09, 1.574449e-10, -2.7336e-10, 1.669792e-08, 
    3.568941e-10, 8.293227e-10, -1.203375e-09, 9.890407e-09, -2.084537e-09, 
    5.398448e-09, 4.162644e-09, 5.255131e-09, 6.374563e-10, -1.520539e-09, 
    -4.036913e-10, -4.187548e-10, 2.579839e-10, 7.018744e-09, -2.768502e-10, 
    -7.111289e-10, -1.147811e-10, 3.399148e-08, 6.756068e-10, 6.079611e-09, 
    -5.284878e-09, -1.272241e-09, -2.30105e-09, -1.290914e-09, -7.511875e-09, 
    -3.405586e-09, 7.932499e-10, -4.044978e-09, 3.323095e-09, 2.004487e-08, 
    4.557194e-09, -1.707974e-09, 2.262746e-08, 4.846754e-10, -4.940262e-10, 
    -4.574739e-09, 2.414708e-10, -3.889511e-11, -2.933227e-09, 6.212232e-10, 
    1.693309e-09, -1.652964e-09, -7.647478e-09, 2.028457e-09, -2.400952e-09, 
    6.51454e-10, -3.289244e-10, 2.435286e-09, -2.227409e-10, -1.155386e-09, 
    -1.911332e-09, 3.198011e-10, 1.170782e-08, -2.707381e-10, -9.832368e-09, 
    1.048704e-09, 1.10104e-09, -5.867037e-10, 5.429968e-09, -4.794174e-10, 
    -2.560228e-11, 3.926402e-09, 5.223857e-10, 2.644818e-11, 3.005596e-10, 
    -1.017099e-09, -4.706635e-11, -6.378968e-10, 1.032845e-10, -1.154802e-09, 
    9.060415e-09, 1.212763e-08, -2.251824e-09, -4.599229e-09, -2.819377e-09, 
    -6.297114e-10, -5.225047e-11, -2.845546e-10, 9.060308e-11, -9.067236e-11, 
    -2.171134e-10,
  -2.66715e-09, 1.078149e-09, 3.821526e-09, 2.113723e-09, -1.637034e-09, 
    1.287788e-09, -9.287533e-09, 1.162277e-09, 4.403944e-09, 1.443652e-09, 
    3.231719e-09, 1.097914e-08, 7.079848e-10, 3.743935e-09, 2.621846e-09, 
    -2.968881e-09, -2.559659e-09, -2.35076e-09, 6.87379e-10, 1.006646e-08, 
    -3.527305e-09, -1.386752e-09, -9.154064e-10, -1.171372e-09, 
    -1.444846e-09, 1.532419e-08, -2.826255e-10, 5.826109e-09, 2.068083e-08, 
    -1.989372e-08, -1.231729e-08, 5.497782e-09, 3.823857e-10, -3.099558e-09, 
    -1.76118e-09, 2.112756e-09, -7.568758e-10, -2.932836e-10, 1.915134e-08, 
    1.19686e-09, 7.267204e-10, -1.600768e-09, 1.178329e-08, -3.288414e-09, 
    3.192326e-09, 7.903679e-09, 1.03677e-08, 7.294005e-10, -2.936804e-09, 
    -4.857661e-10, 1.957545e-11, 1.283013e-09, 1.153921e-08, -7.480707e-10, 
    2.239318e-10, -7.531753e-11, 3.989021e-08, 8.432665e-10, 3.018923e-08, 
    -9.280505e-09, -6.142102e-09, -1.58991e-09, -1.525052e-09, -9.701011e-10, 
    -1.549586e-09, 9.378994e-09, -1.706326e-09, 1.157309e-08, 2.216484e-08, 
    3.615128e-09, -1.029946e-09, 9.409803e-09, 2.465299e-10, 7.433414e-10, 
    -6.75294e-10, 2.150387e-10, -1.937437e-10, -4.068497e-09, 9.085639e-10, 
    4.305662e-09, -1.226226e-09, -1.123948e-08, 1.838032e-09, 5.156835e-10, 
    -2.538513e-09, 3.019409e-09, 1.600938e-09, -3.017249e-10, -1.404328e-09, 
    -2.554231e-09, 8.950906e-09, 1.884126e-08, -1.104397e-09, -2.297648e-08, 
    3.126388e-11, 2.032164e-09, -7.254812e-10, 3.092907e-09, -6.148753e-10, 
    -2.141405e-10, 3.064429e-09, -2.273325e-09, 1.90532e-10, 1.490825e-10, 
    -6.928076e-10, -2.078764e-10, 3.290666e-10, 2.527941e-09, -1.289038e-09, 
    7.837116e-09, 5.006541e-09, -1.349179e-09, -6.77943e-09, -2.851834e-09, 
    2.860929e-10, -6.667733e-11, -1.491856e-10, 9.781509e-11, -9.81828e-11, 
    3.432206e-10,
  -1.217586e-09, 3.70278e-10, -1.776584e-09, -9.907808e-10, -1.461558e-09, 
    -1.784713e-09, -1.237316e-08, 2.385718e-10, 4.657181e-09, 2.079332e-10, 
    1.205024e-09, 6.363337e-09, -2.07848e-09, -1.286367e-10, 7.013227e-09, 
    -3.63512e-09, -4.3216e-09, -2.609795e-09, -1.299512e-10, 1.870751e-08, 
    -4.485628e-09, -1.327635e-09, -1.853266e-09, -8.614052e-10, 
    -1.300293e-09, 4.606363e-09, -1.781245e-09, -8.752352e-09, 4.453284e-09, 
    -9.483017e-09, -1.921785e-08, 3.522416e-09, 7.37657e-10, -3.284754e-09, 
    -3.542993e-09, 5.039851e-09, -1.444306e-09, -1.929976e-10, 3.376914e-08, 
    2.002782e-09, 1.637659e-10, -7.057849e-09, 1.599118e-08, -5.055756e-09, 
    9.732673e-09, 1.024841e-08, 1.691666e-08, 1.06229e-09, -4.25232e-09, 
    -5.849508e-10, 8.3336e-10, 3.500645e-09, 1.840112e-08, -1.062517e-09, 
    1.950312e-09, 6.372147e-11, 4.568193e-08, 1.164267e-09, 6.66083e-08, 
    -1.147341e-08, -1.28349e-08, 7.92852e-10, -1.011699e-09, 2.044544e-10, 
    -3.401317e-09, 1.328112e-08, 3.325965e-09, 2.4965e-08, 2.225772e-08, 
    1.100608e-08, -1.245496e-09, 2.560739e-09, -2.601723e-10, 2.092463e-09, 
    3.169964e-09, 1.538751e-10, -4.267946e-10, -6.213384e-09, 1.225072e-09, 
    1.943306e-09, -3.153161e-09, -1.650228e-08, 1.078064e-09, 2.800107e-09, 
    -1.624358e-09, 3.628315e-09, -3.220748e-10, -5.185825e-10, -3.598485e-09, 
    -2.939231e-09, 1.190307e-08, 2.512612e-08, -2.615323e-09, -3.734469e-08, 
    3.820787e-09, 3.248454e-09, -5.36295e-10, -1.580872e-09, -9.949304e-10, 
    -6.467644e-10, 1.104809e-09, -6.137686e-09, 3.541025e-10, 6.282264e-11, 
    -1.896467e-09, -2.184208e-09, -3.353193e-09, -1.071271e-09, 
    -3.608193e-09, 6.66995e-09, 2.325521e-09, -1.000274e-09, -5.694972e-09, 
    -3.017419e-09, 1.222304e-09, -9.993641e-11, -6.211565e-11, 8.468604e-11, 
    -9.34719e-11, -2.208935e-10,
  2.116565e-09, -7.095196e-10, -3.829996e-09, -2.260037e-09, -9.432597e-10, 
    -2.720071e-09, -4.970843e-09, -8.145662e-11, 3.707441e-09, 1.193484e-09, 
    -1.876515e-09, 4.379615e-09, -2.710919e-09, 3.370246e-09, 5.575714e-09, 
    -9.632064e-10, -5.501363e-09, -5.164452e-09, -1.569568e-09, 2.75428e-08, 
    1.41614e-09, -2.299885e-09, -1.299611e-09, 2.345928e-10, -5.261427e-10, 
    1.691433e-09, 3.990465e-09, -1.815005e-08, -1.301885e-09, -2.96086e-09, 
    -1.930027e-08, -1.007948e-09, 1.779995e-09, -5.295647e-09, -3.196078e-09, 
    5.837137e-09, -1.465361e-09, -1.491074e-10, 6.257829e-08, 2.044686e-09, 
    -4.617618e-10, -1.112335e-08, 1.718109e-08, -6.531527e-09, 3.083875e-08, 
    -6.669552e-09, 1.837807e-08, 6.110184e-09, -6.505944e-09, -8.865157e-10, 
    2.302443e-09, 3.115701e-09, 2.680973e-08, -6.043592e-10, 4.259228e-09, 
    2.409308e-10, 5.23554e-08, 1.727636e-09, 8.471736e-08, -9.675233e-09, 
    -9.472274e-09, 4.08528e-09, -2.913225e-10, -1.295018e-09, -4.886249e-09, 
    -4.390984e-09, 1.047499e-08, 6.568519e-08, 2.777421e-08, 2.025195e-08, 
    -2.01311e-09, 1.797406e-08, -2.290221e-10, 1.765784e-09, 7.703687e-09, 
    1.932676e-12, -5.889831e-10, -9.2856e-09, 1.670074e-09, -4.88285e-10, 
    -4.826461e-09, -2.315576e-08, 2.813749e-12, -8.249685e-10, 2.424997e-09, 
    3.397986e-09, -3.473701e-09, -6.508003e-10, -4.786394e-09, -1.764818e-09, 
    9.442715e-09, 2.949646e-08, -3.269022e-09, -3.536687e-08, 5.232948e-09, 
    4.390637e-09, 1.522267e-11, -1.071641e-08, -1.164949e-09, -1.287879e-09, 
    9.227961e-10, 4.429271e-09, 2.279563e-10, 1.670024e-10, -6.57684e-09, 
    -1.746798e-10, 1.381522e-09, -1.252624e-08, -3.627918e-09, 8.176357e-09, 
    3.053401e-09, -1.410456e-09, -1.735316e-09, -3.752689e-09, -1.603837e-09, 
    -1.602189e-10, 2.217106e-10, 1.061835e-10, -5.16529e-11, -1.063881e-09,
  4.074593e-09, -4.077549e-09, -3.462048e-09, -1.448541e-09, -4.687308e-10, 
    -1.297508e-09, 2.563979e-09, -1.625324e-09, 4.259107e-09, 2.816137e-09, 
    -3.557091e-09, 2.215756e-10, -4.941342e-09, 9.965788e-10, 6.11692e-09, 
    -6.478444e-10, -8.387724e-09, -5.702759e-09, -2.680224e-09, 2.823566e-08, 
    5.27848e-09, -6.878338e-09, 1.105263e-09, 2.890886e-09, -5.915695e-10, 
    8.771508e-10, 2.1034e-08, -2.39898e-08, 1.464986e-08, 4.110802e-09, 
    -1.863162e-08, -5.283539e-09, 7.484573e-10, -9.29731e-09, -1.847923e-09, 
    5.83475e-09, -3.433035e-09, -6.834e-11, 9.243729e-08, 8.022027e-10, 
    -1.228e-09, -1.750777e-10, 1.684168e-08, -7.956506e-09, 6.742408e-08, 
    -2.565042e-08, 1.788763e-08, 1.209891e-08, -9.033704e-09, -1.247439e-09, 
    6.019704e-09, -1.116632e-09, 3.770327e-08, -5.158199e-10, 7.989904e-09, 
    4.327205e-10, 6.098128e-08, 2.344296e-09, 7.301919e-08, -2.489998e-09, 
    5.320544e-11, 5.816844e-09, 4.919229e-10, -3.693333e-09, -8.352732e-09, 
    -9.169582e-09, 2.238573e-08, 7.652574e-08, 2.907319e-08, 2.332882e-08, 
    -1.667502e-09, 2.270468e-08, -5.8605e-09, -3.249738e-10, 1.265342e-08, 
    -1.969056e-10, -8.225953e-10, -1.292986e-08, 2.174991e-09, 1.580793e-08, 
    -4.035229e-09, -3.490874e-08, -6.886012e-10, 5.447873e-10, 7.089e-09, 
    1.97798e-09, -4.100229e-09, -1.654541e-09, -1.107539e-08, -1.564757e-09, 
    2.376737e-09, 3.208093e-08, -1.427537e-09, 1.181083e-08, 6.488676e-09, 
    5.420162e-09, 3.139121e-10, -1.048409e-08, -1.370609e-09, -2.097022e-09, 
    2.623324e-10, 1.544042e-08, -3.227321e-10, 4.61327e-10, -2.034653e-09, 
    3.323407e-09, 1.361116e-09, -1.989628e-08, 7.01715e-09, 1.191142e-08, 
    4.07266e-09, -5.932975e-09, 1.246178e-09, -4.986077e-09, -8.025211e-09, 
    -2.664819e-10, 7.61105e-10, 1.443041e-10, 2.00906e-11, -1.520561e-09,
  5.157005e-09, -6.970311e-09, -2.581203e-09, -8.948859e-10, -6.651248e-10, 
    1.754756e-09, 4.868639e-09, -1.245297e-08, 4.961123e-09, 1.693479e-09, 
    -7.656809e-10, -2.753382e-09, -2.899299e-09, -4.272522e-09, 1.253102e-08, 
    1.408084e-09, -1.309055e-08, -3.424418e-09, -3.373181e-09, 2.312601e-08, 
    -1.129933e-09, -1.889049e-08, 2.191769e-09, 4.16162e-09, -4.774847e-12, 
    1.415401e-11, 8.169297e-08, -1.582839e-08, 6.334631e-09, 1.524359e-08, 
    -2.030998e-08, -6.204004e-09, -2.967681e-09, -1.61545e-08, 9.815722e-10, 
    4.070785e-09, -4.729259e-09, 1.698623e-10, 1.090967e-07, -2.165887e-09, 
    -2.726131e-09, 6.957805e-09, 1.800909e-08, -1.005904e-08, 8.417152e-08, 
    -1.106849e-08, 1.682685e-08, 1.539942e-08, -8.146289e-09, -1.688331e-09, 
    7.747452e-09, -8.493714e-09, 5.277012e-08, -8.58131e-10, 1.466732e-08, 
    5.491358e-10, 6.702766e-08, -4.265757e-10, 4.617982e-08, -1.852598e-09, 
    -4.142237e-09, 5.143306e-09, 1.965759e-09, -4.27384e-09, -9.097141e-09, 
    -2.344933e-08, 3.496285e-08, 7.204687e-08, 3.740644e-08, 1.263055e-08, 
    -3.050332e-09, 2.204939e-08, -2.643316e-08, -2.060005e-10, 1.407334e-08, 
    -4.561684e-10, -8.275407e-10, -1.474524e-08, 2.301164e-09, 2.61781e-08, 
    -4.824983e-09, -4.283214e-08, -1.189619e-09, 9.183054e-10, -1.706837e-09, 
    9.183054e-10, -2.740308e-09, -1.988781e-09, -1.077711e-08, -2.270895e-09, 
    4.374101e-10, 3.411404e-08, 6.288587e-10, 7.846256e-08, 6.207244e-09, 
    6.480229e-09, -1.683452e-09, -7.013909e-09, -4.95163e-10, -3.068419e-09, 
    -2.785328e-10, 7.383381e-09, -9.144543e-10, 3.878355e-10, 1.070981e-08, 
    2.151864e-09, -1.189125e-08, 1.605997e-09, 2.066719e-08, 9.769053e-09, 
    1.959165e-09, -1.015371e-08, 3.821526e-09, -5.887728e-09, -1.270809e-08, 
    -3.471655e-10, 1.212292e-09, 1.930474e-10, 7.223733e-11, -1.192291e-09,
  5.740503e-09, -4.38547e-09, -4.413835e-09, -4.747335e-09, -1.180467e-09, 
    2.404363e-09, 2.832962e-09, -2.894546e-08, 2.447223e-09, -7.679546e-10, 
    -9.75092e-10, -3.361777e-09, 9.043788e-10, -4.907633e-09, 1.211055e-08, 
    1.460677e-09, -1.832848e-08, -2.32734e-09, -2.468084e-09, 2.056839e-08, 
    -2.36065e-09, -7.807444e-10, -7.58962e-09, 5.325376e-09, 7.485141e-10, 
    -2.978027e-10, 9.444301e-08, 7.728488e-09, 1.776554e-07, 3.292655e-09, 
    -1.748396e-08, -7.800395e-09, -9.802136e-09, -2.695487e-08, 8.698748e-10, 
    1.207241e-09, -7.856317e-09, 5.946035e-10, 1.055755e-07, -6.05403e-09, 
    -8.171992e-09, 7.742642e-09, 1.945041e-08, -1.065912e-08, 7.019491e-08, 
    1.584948e-08, 1.476693e-08, 1.472706e-08, 2.760647e-09, -2.287322e-09, 
    6.653991e-09, -8.069094e-09, 7.295377e-08, -1.950832e-09, 2.23098e-08, 
    5.209415e-10, 6.503024e-08, -6.385028e-09, 2.139267e-08, -3.754934e-09, 
    -7.246115e-09, 4.501771e-09, 3.893376e-09, -4.881383e-09, -1.199685e-08, 
    -4.66847e-08, 2.515981e-08, 7.482544e-08, 4.028038e-08, -8.256563e-09, 
    -2.493266e-09, 8.715176e-09, -1.878584e-08, -1.750323e-09, 1.144078e-08, 
    -8.171241e-10, -9.615775e-10, -1.520225e-08, 1.408273e-09, 2.081191e-08, 
    -8.139693e-09, -5.271766e-08, -2.185175e-09, 7.790959e-10, -4.614947e-09, 
    -3.592504e-11, -4.132971e-09, 2.665956e-11, -4.224752e-09, -6.424472e-09, 
    -7.275958e-11, 3.57524e-08, 2.759251e-09, 1.462991e-07, 5.625054e-09, 
    8.262259e-09, -8.843881e-09, 1.440191e-08, 1.444903e-09, -3.916034e-09, 
    -1.103729e-09, -1.153932e-09, -1.814836e-09, -9.940493e-11, 4.817082e-09, 
    -3.897696e-09, -7.785445e-09, 1.826908e-08, 1.724572e-08, 3.17732e-09, 
    -1.079172e-09, -7.169831e-09, 2.318245e-09, -5.921265e-09, -2.029321e-08, 
    -5.108348e-10, 1.72389e-09, 2.79627e-10, 1.016183e-10, 1.558078e-09,
  3.238938e-09, -1.408239e-09, -4.328456e-09, -1.88154e-08, -2.962679e-10, 
    2.486388e-09, -2.751221e-10, -2.876351e-08, -1.510955e-09, -7.729739e-09, 
    -2.928289e-09, 6.946834e-10, 8.184884e-10, -1.893909e-09, -1.586102e-09, 
    2.614808e-09, -2.049576e-08, 8.477059e-10, -4.304916e-09, 1.934626e-08, 
    -5.643017e-09, 6.687571e-09, -1.369472e-08, -3.902301e-10, 1.501576e-09, 
    -5.603056e-10, 6.708598e-08, 1.544731e-08, 8.523955e-09, -1.716808e-08, 
    -7.152209e-09, -2.245542e-09, 7.789367e-09, -2.922172e-08, -3.039588e-09, 
    2.455636e-11, -8.739898e-09, 1.348155e-09, 1.09752e-07, -1.013713e-08, 
    -2.331588e-08, 3.53964e-09, 1.819112e-08, -1.120574e-08, 5.803122e-08, 
    2.407307e-08, 1.436712e-08, 1.474244e-08, 2.863567e-08, -3.198494e-09, 
    3.709779e-09, -3.095067e-09, 9.930095e-08, -9.977155e-11, 3.171948e-08, 
    3.78094e-10, 5.89759e-08, -8.73614e-09, 1.093903e-08, -1.395676e-08, 
    1.446926e-08, 6.283756e-09, 2.953868e-09, -6.666096e-09, -1.878127e-08, 
    -5.447532e-08, 1.645634e-08, 6.573504e-08, 4.15933e-08, -1.086005e-08, 
    -4.599769e-09, -1.677228e-08, -1.496323e-08, -5.037066e-09, 1.161241e-08, 
    -1.312856e-09, -1.356803e-09, -7.88161e-09, -4.141398e-10, 4.58914e-09, 
    -7.990195e-09, -8.475634e-08, -3.323493e-09, 1.36771e-09, -2.491902e-09, 
    -7.323536e-09, -4.138883e-09, 3.94482e-09, -1.204418e-09, -5.304344e-09, 
    -1.778403e-09, 3.019682e-08, 3.904773e-09, 1.67003e-07, 4.734488e-09, 
    1.071627e-08, -1.833332e-08, 5.045263e-08, 4.157357e-09, -4.285016e-09, 
    -1.162618e-09, -9.692123e-10, -5.962054e-09, -6.72248e-10, -8.692325e-09, 
    -5.347317e-09, -3.833009e-09, 6.700077e-09, 5.230788e-09, 1.532499e-10, 
    -4.681056e-09, -3.470859e-10, 3.012701e-12, -4.931564e-09, -2.261174e-08, 
    -7.871904e-10, 2.224667e-09, 3.989289e-10, 9.428547e-11, 5.397283e-09,
  -9.496262e-10, -1.720991e-09, 4.769163e-10, -3.845162e-08, -7.074163e-10, 
    5.199468e-09, 6.355094e-11, -9.516611e-09, -1.973154e-08, -1.134907e-08, 
    -1.239528e-09, 6.299445e-09, 1.663238e-10, 2.993943e-10, -6.27108e-09, 
    6.165507e-09, -2.276552e-08, 5.881105e-09, -8.725856e-09, 1.538069e-08, 
    1.085147e-08, 2.684203e-09, -1.03114e-10, -8.589041e-09, 2.516799e-09, 
    -1.006129e-09, 1.905107e-08, 1.524614e-08, -1.925018e-07, -3.862363e-08, 
    7.358665e-09, 2.927095e-09, -4.438562e-09, -9.70374e-10, -1.395711e-08, 
    1.382205e-09, -5.628255e-09, 2.308553e-09, 1.682106e-07, -1.494915e-08, 
    -4.160231e-08, 5.450488e-09, 1.585664e-08, -1.249979e-08, 2.875333e-08, 
    -5.896936e-10, 1.968019e-08, 5.922843e-09, 3.80813e-08, -4.274494e-09, 
    -4.230074e-10, -4.120238e-09, 1.259579e-07, 3.290325e-10, 3.77268e-08, 
    1.944329e-10, 6.67207e-08, -8.153962e-10, 1.161701e-08, -2.919738e-08, 
    2.138808e-08, 6.10089e-09, 2.059835e-09, -9.268138e-09, -2.297523e-08, 
    -1.292887e-08, 1.121168e-08, 4.631346e-08, 3.240979e-08, -9.56652e-09, 
    -2.697163e-08, -5.248421e-08, -9.164637e-09, -5.682466e-09, 2.803836e-08, 
    -1.864578e-09, -2.65338e-10, 1.844469e-09, -3.052296e-09, -4.208118e-10, 
    -5.193414e-09, -1.213862e-07, -5.302184e-09, -3.482796e-10, 
    -1.076899e-09, -1.657588e-08, -2.624802e-09, 5.971458e-09, -1.392445e-08, 
    1.138565e-08, -3.609557e-09, 2.588591e-08, 3.833094e-09, 1.268312e-07, 
    -1.725823e-09, 1.174726e-08, -2.140051e-08, 9.434405e-08, 5.515346e-09, 
    -5.156392e-09, -7.800054e-10, 1.469175e-09, -6.23341e-09, -2.531159e-09, 
    -1.824844e-08, -4.668266e-09, -1.548204e-08, -2.339777e-08, 1.021931e-09, 
    -3.744333e-09, -9.6245e-09, 1.909484e-09, -1.382659e-09, -4.567369e-09, 
    -4.30839e-09, -1.146043e-09, 2.524835e-09, 4.393286e-10, 5.907452e-11, 
    7.865026e-09,
  -3.967784e-09, -1.827516e-09, 1.565161e-08, -3.284379e-08, -2.403226e-09, 
    9.363248e-09, -5.373977e-10, 7.81904e-09, -3.24186e-08, -7.027438e-09, 
    1.848321e-09, 7.463655e-09, -9.796395e-10, 1.009016e-08, -1.909939e-10, 
    4.839102e-09, -3.085611e-08, 9.67583e-09, -4.898965e-09, 6.361347e-09, 
    5.363529e-08, -2.381285e-08, -9.925884e-09, -2.065462e-09, 1.790681e-09, 
    -7.046765e-09, 1.327862e-09, 1.076103e-08, -1.53348e-07, -5.749507e-08, 
    7.996346e-08, 2.00024e-08, 2.636421e-08, 3.906871e-08, -2.221043e-08, 
    1.969579e-08, -1.25284e-09, 3.675225e-09, 9.30396e-08, -5.613094e-08, 
    -5.278248e-08, 5.916263e-09, 1.777215e-08, -1.084746e-08, -6.616006e-09, 
    -3.216837e-08, 3.117015e-08, -3.484101e-08, 4.633062e-08, -5.22148e-09, 
    -5.943178e-09, -2.214847e-08, 1.461221e-07, -4.086973e-09, 4.402902e-08, 
    -2.65004e-10, 6.566052e-08, -3.374271e-09, 7.79554e-09, -1.844734e-08, 
    4.323738e-09, 2.605134e-09, 1.956437e-09, -8.32606e-09, -2.275542e-08, 
    6.315076e-09, 2.251094e-07, 2.656054e-08, 2.143861e-08, 1.192927e-08, 
    -1.281796e-08, -1.317649e-07, -1.176227e-08, -1.185413e-09, 5.276977e-08, 
    -2.23406e-09, 1.124263e-09, 2.442945e-08, -5.781976e-09, -1.210879e-09, 
    -3.961361e-09, -1.367959e-07, -6.574396e-09, -4.860226e-09, 1.09718e-08, 
    1.947808e-08, 3.326477e-10, 4.835329e-09, -4.048414e-08, 3.233527e-08, 
    -3.513151e-09, 2.973113e-08, 3.636245e-09, 5.582102e-08, -1.018964e-08, 
    8.796564e-09, -1.54092e-08, 3.842626e-08, 4.859544e-09, -8.199549e-09, 
    3.763034e-11, -1.548116e-09, 1.455255e-09, -8.530037e-09, -2.299612e-08, 
    -7.022095e-09, -2.740092e-08, -4.000538e-08, -1.655508e-09, 
    -3.620016e-09, -1.099647e-08, 4.398544e-10, -8.345751e-10, -4.042022e-09, 
    8.807206e-09, -1.369074e-09, 2.784859e-09, 3.049543e-10, 1.774936e-11, 
    3.272021e-09,
  3.833446e-08, 3.94067e-09, 2.980636e-08, 4.162933e-08, 2.377135e-09, 
    1.137965e-08, 1.396643e-10, 1.212157e-08, -1.934023e-08, 3.000139e-09, 
    5.265804e-09, 4.898936e-09, -7.538006e-10, 2.365863e-08, 2.647255e-09, 
    2.025352e-09, -4.621435e-08, 1.906238e-08, 6.489145e-09, 4.537867e-09, 
    7.182251e-08, -1.892676e-08, -4.790371e-08, -3.043425e-08, -1.723396e-08, 
    -9.390931e-09, -9.959848e-08, 7.86298e-09, -1.265524e-07, -7.024875e-08, 
    2.127525e-07, 1.518085e-07, 3.45853e-08, 1.076331e-07, -4.094858e-08, 
    5.821386e-08, 5.321295e-09, 6.576101e-09, 1.276663e-08, -6.10365e-08, 
    -6.618435e-08, 4.503306e-09, 1.851868e-08, -1.053642e-08, -1.618224e-08, 
    -1.010011e-07, 3.972013e-08, -8.655934e-08, 4.934585e-08, -6.080803e-09, 
    -1.258833e-08, -4.921236e-08, 1.37078e-07, -9.812777e-09, 4.733673e-08, 
    -1.431715e-09, 3.122449e-08, -1.937489e-08, -2.176648e-10, 2.487582e-09, 
    2.593765e-10, 4.710614e-10, 2.012996e-09, -5.024695e-09, -3.061085e-08, 
    5.948948e-09, 2.075764e-07, 1.707195e-08, 1.919472e-08, 2.905e-08, 
    6.790685e-09, -1.674298e-07, -2.07794e-08, -1.817341e-09, 5.566238e-08, 
    -3.6556e-10, 2.521929e-09, 4.496576e-08, -8.5587e-09, 2.116843e-08, 
    -2.181082e-09, -1.320024e-07, -7.71297e-09, -8.769291e-09, 1.325867e-08, 
    2.431765e-07, 5.714071e-09, 3.444086e-09, -5.946942e-08, 5.716248e-08, 
    -1.815295e-09, 3.113697e-08, 2.540048e-09, 4.987328e-09, -7.55719e-08, 
    1.881744e-10, -4.702463e-09, 4.00932e-08, 1.765613e-09, -1.298068e-08, 
    5.974243e-11, -5.443404e-09, 4.878537e-09, -1.338243e-08, -7.294938e-08, 
    -5.410072e-09, -4.163081e-08, -5.805902e-08, -5.117897e-09, 9.385417e-10, 
    -7.453366e-09, -3.134062e-09, -3.912533e-10, -1.641467e-09, 1.689898e-09, 
    -1.602052e-09, 3.621807e-09, 9.573498e-11, -4.445155e-11, -9.07761e-09,
  1.035703e-07, 7.846552e-09, 3.42086e-08, 1.57124e-07, 2.185971e-08, 
    1.602268e-08, 6.22174e-09, 1.102342e-08, 9.911446e-09, 4.603294e-09, 
    4.209255e-09, 1.454168e-09, -2.130946e-09, 2.621414e-08, 4.592948e-09, 
    -4.380659e-09, -5.089855e-08, 3.41272e-08, -6.264277e-08, 1.354704e-08, 
    4.375966e-08, -1.422188e-08, -3.567948e-09, -3.559228e-08, -1.095759e-08, 
    1.725198e-09, -5.717457e-07, 2.376282e-09, -9.026235e-08, -7.360484e-08, 
    1.03009e-07, 2.017429e-07, -7.629717e-08, 1.031656e-07, -8.241102e-08, 
    8.56827e-08, 1.58022e-08, 9.792686e-09, 3.232549e-08, -5.818332e-08, 
    -8.700181e-08, 2.445404e-09, 1.284081e-08, -1.414258e-08, -1.343824e-08, 
    -1.705847e-07, 4.864756e-08, -1.321069e-07, 4.696274e-08, -6.338354e-09, 
    -1.916291e-08, -5.301138e-08, 9.96698e-08, -9.877226e-09, 4.702463e-08, 
    -2.292097e-09, 1.297121e-08, -3.217912e-08, 4.415415e-09, 2.949196e-08, 
    2.16744e-09, 1.170974e-11, -1.017611e-09, -1.793389e-09, -5.331751e-08, 
    -7.098492e-09, 6.638334e-08, 2.101115e-08, 2.05581e-08, 3.923844e-08, 
    -6.288474e-09, -1.028878e-07, -3.072444e-08, -3.023729e-09, 3.792193e-08, 
    1.726107e-09, 3.224386e-09, 7.076528e-08, -1.064311e-08, 3.276774e-07, 
    1.965077e-10, -1.401269e-07, -1.466867e-08, -7.71729e-09, 1.893568e-09, 
    1.973376e-07, 2.363436e-09, 6.942855e-10, -7.466586e-08, 5.980939e-08, 
    -4.445155e-11, 2.105139e-08, 2.695373e-09, -4.027108e-08, -5.885693e-08, 
    -1.312969e-08, 1.519738e-08, 7.6883e-08, 4.082494e-09, -1.710439e-08, 
    -6.32906e-09, -5.120881e-11, 3.297657e-09, -1.704469e-08, -9.504572e-08, 
    -1.041337e-08, -5.449567e-08, -5.886477e-08, -9.944529e-09, 3.85171e-10, 
    2.516799e-09, -3.52793e-09, -2.285105e-09, 9.716814e-10, -3.098648e-09, 
    -1.908825e-09, 4.984997e-09, -3.472174e-10, -1.080878e-10, -1.119997e-08,
  1.692273e-07, 5.966683e-09, 1.982579e-08, 1.545648e-07, 1.328266e-08, 
    1.881216e-08, 2.321832e-08, 7.107133e-10, 3.211375e-08, 5.2475e-09, 
    3.564082e-11, -2.031868e-09, -1.510159e-09, -3.131504e-10, 1.941811e-08, 
    -1.246721e-08, -6.16284e-08, 4.759482e-08, -1.536782e-07, 2.19357e-08, 
    7.60366e-09, -1.476963e-09, 2.250482e-08, 1.798986e-08, 7.68847e-09, 
    6.357652e-09, -4.370272e-07, 5.314007e-09, -9.332456e-08, -7.951229e-08, 
    -1.428174e-08, 7.284126e-08, -5.775365e-08, 5.344106e-08, -1.120902e-07, 
    8.910439e-08, 2.503506e-08, 1.255344e-08, 7.796024e-08, -3.435912e-08, 
    -1.115385e-07, 1.946717e-09, 9.416482e-09, -1.973755e-08, -1.316829e-08, 
    -1.918353e-07, 6.545196e-08, -1.399086e-07, 3.551623e-08, -6.412407e-09, 
    -2.766764e-08, -4.573002e-08, 5.023142e-08, -5.302388e-09, 5.19153e-08, 
    -1.789147e-09, 1.353914e-08, -9.027124e-08, 1.597354e-08, 4.290735e-08, 
    2.11287e-10, 1.705303e-13, 2.57366e-08, -6.287259e-09, -5.968305e-08, 
    -2.930204e-08, 1.132088e-08, 2.042287e-08, 1.972506e-08, 4.629027e-08, 
    2.261896e-08, -1.342159e-07, -2.602343e-08, -1.03492e-08, 3.204543e-08, 
    -1.029974e-08, 1.989363e-09, 8.337108e-08, -1.180531e-08, 2.923915e-07, 
    2.669765e-09, -1.547256e-07, -2.820423e-08, -5.793311e-09, -9.334315e-09, 
    -1.054362e-07, -1.484031e-07, 7.947108e-09, -9.637376e-08, 5.26033e-08, 
    -5.200604e-10, 1.260222e-08, 3.908156e-09, -8.943837e-08, -2.335298e-09, 
    -2.528021e-08, 5.654903e-08, 5.818487e-08, 9.078065e-09, -2.021076e-08, 
    -2.36634e-08, 1.026951e-08, 1.337905e-08, -1.686367e-08, -4.753537e-08, 
    -4.415045e-08, -4.539953e-08, -5.425562e-08, -1.129609e-08, 
    -2.057448e-09, 1.274447e-08, 1.096453e-09, -2.159993e-09, -4.152241e-09, 
    -3.769117e-09, -1.980538e-09, 6.89073e-09, -6.206804e-10, -1.836398e-10, 
    5.392224e-09,
  1.594543e-07, 1.952742e-09, 2.308809e-09, 4.771795e-08, 6.602875e-09, 
    1.816835e-08, 4.092732e-08, -1.415009e-08, 1.13443e-08, 2.532545e-09, 
    4.100116e-10, -2.111676e-09, -2.955687e-09, -2.611301e-08, 2.26392e-08, 
    -1.385666e-08, -7.303769e-08, 6.360119e-08, -1.323935e-07, 2.863879e-08, 
    -2.132373e-08, 1.93296e-09, 1.016389e-08, 7.630263e-09, 1.055145e-08, 
    1.047624e-10, -6.845443e-08, 7.67767e-09, -8.683145e-08, -1.062454e-07, 
    -1.446944e-08, 2.566424e-09, 2.751568e-08, 4.922055e-08, -1.210164e-07, 
    8.573107e-08, 2.835333e-08, 1.53078e-08, 1.207122e-07, 3.47755e-08, 
    -7.550076e-08, 7.067172e-09, 7.549573e-09, -2.661516e-08, -2.066434e-08, 
    -1.62342e-07, 9.297935e-08, -9.804316e-08, 1.604568e-08, -6.921532e-09, 
    -3.024094e-08, -3.471888e-08, 1.412011e-08, -2.572404e-09, 5.88093e-08, 
    -3.529976e-09, 3.744901e-09, -4.467476e-08, 2.402589e-08, 5.671765e-08, 
    -2.766853e-09, -5.886136e-10, 9.73651e-08, -1.550023e-08, -3.794447e-08, 
    -4.080295e-08, -1.78249e-08, 3.454949e-08, 1.690904e-08, 3.649023e-08, 
    -1.061778e-09, -3.513327e-08, -8.157997e-09, -9.71778e-09, 5.935705e-08, 
    -2.700796e-08, -9.557084e-10, 8.531879e-08, -1.206201e-08, 2.416385e-08, 
    2.61997e-09, -1.682859e-07, -2.672567e-08, -6.106688e-10, -9.694475e-09, 
    2.976498e-08, -3.435691e-07, 2.070971e-08, -1.358998e-07, 3.826983e-08, 
    3.628315e-10, 6.463517e-09, 3.627349e-09, -1.542383e-07, 1.126449e-08, 
    -3.000955e-08, 5.465048e-08, 5.302525e-09, 1.626057e-08, -2.367705e-08, 
    -4.01472e-08, 6.90531e-09, 1.105038e-08, -1.180918e-08, -2.30205e-08, 
    -5.36358e-08, -2.778819e-08, -3.771362e-08, -5.642448e-09, -3.323692e-09, 
    7.880487e-09, -5.246079e-10, -5.794334e-09, -2.138239e-08, -3.038565e-09, 
    -1.806461e-09, 9.458958e-09, -6.052048e-10, -2.798402e-10, 4.353353e-09,
  6.004416e-08, 2.606839e-10, -1.298122e-08, -2.641264e-08, 8.193524e-09, 
    1.500769e-08, 4.764013e-08, -1.984529e-08, -1.299088e-08, -6.327014e-09, 
    -3.366949e-09, 9.958967e-11, -6.706387e-10, -1.35833e-09, 1.554724e-08, 
    -9.282463e-09, -8.518853e-08, 5.928621e-08, -2.408994e-08, 2.518266e-08, 
    -2.458773e-08, 1.031594e-09, 5.594529e-10, -2.594675e-09, 9.346195e-10, 
    -2.70154e-08, -3.91118e-08, 1.385206e-08, -8.060363e-08, -1.611298e-07, 
    1.054809e-08, -3.581022e-08, 5.013055e-08, 6.511414e-08, -1.402152e-07, 
    7.541928e-08, 2.34708e-08, 1.803672e-08, 1.198259e-07, 1.122698e-07, 
    1.991493e-08, 6.934329e-09, 9.30811e-09, -3.053308e-08, 3.737796e-09, 
    -1.266612e-07, 1.312293e-07, 1.574787e-08, -2.026636e-08, -9.11308e-09, 
    -2.807656e-08, -3.474827e-08, -1.659579e-08, -9.020369e-10, 5.929571e-08, 
    -1.787726e-09, -7.367476e-09, -3.960334e-08, 3.623516e-08, 7.095881e-08, 
    -2.387196e-09, -5.418201e-09, 1.144729e-07, -3.278381e-08, -2.545696e-08, 
    -2.364084e-08, -4.243213e-08, 3.929017e-08, 1.616445e-08, 3.243156e-08, 
    -4.283916e-07, -1.277317e-08, 8.79254e-10, 7.42682e-09, 7.363774e-08, 
    -2.916227e-08, -3.688839e-09, 7.26877e-08, -1.196953e-08, 1.697242e-08, 
    6.666312e-09, -1.371798e-07, -2.030163e-09, -4.887966e-09, -4.732783e-10, 
    1.075647e-07, -1.412068e-07, 2.859576e-08, -1.609892e-07, 3.152758e-08, 
    -1.087494e-08, -4.730378e-08, 1.100261e-09, -1.581744e-07, 1.559215e-09, 
    -1.679049e-08, -1.796912e-09, 1.39745e-08, 6.130108e-09, -2.65914e-08, 
    -1.914805e-08, -1.465712e-08, 5.719457e-09, -4.43373e-09, -3.426999e-08, 
    -3.836806e-08, -4.381866e-08, -2.383706e-08, 4.970047e-09, 5.842139e-09, 
    -2.444267e-11, -4.874209e-09, -1.45269e-08, -4.262472e-08, -1.173362e-09, 
    -1.662352e-09, 1.116909e-08, -9.724381e-10, -3.651408e-10, -7.855624e-08,
  3.147119e-08, -7.88134e-10, -2.689188e-08, -3.356621e-08, 1.59402e-08, 
    2.361702e-08, 5.438113e-08, -1.949633e-08, -3.572762e-08, 9.386554e-10, 
    -1.203375e-10, -7.030962e-10, -4.512515e-09, 3.48831e-09, 1.679354e-08, 
    -7.621669e-09, -8.421129e-08, 3.185858e-08, 1.27153e-08, -2.361105e-09, 
    -1.021823e-08, -2.419824e-10, 3.123546e-10, -1.500268e-09, -1.832234e-09, 
    -1.220539e-07, -2.663086e-08, 2.779365e-08, -7.317379e-08, -1.820461e-07, 
    4.851591e-08, -5.587088e-08, 3.829274e-08, 8.441367e-08, -1.447324e-07, 
    4.215968e-08, 1.789271e-08, 2.038006e-08, 1.153962e-07, 1.844324e-07, 
    6.340102e-08, 4.367223e-09, 1.399542e-08, -3.087489e-08, 3.435929e-08, 
    -1.221771e-07, 1.762832e-07, 1.488115e-07, -6.040631e-08, -1.092037e-08, 
    -2.303119e-08, -4.027669e-08, -3.677433e-08, -8.375424e-10, 5.447305e-08, 
    -1.697572e-09, 2.236101e-08, -2.804312e-10, 5.827022e-08, 6.751451e-08, 
    2.01851e-10, -7.347069e-09, 1.59611e-07, -3.241879e-08, -4.539121e-08, 
    1.888736e-09, -1.541423e-09, 3.800739e-08, 1.692621e-08, 2.957228e-08, 
    -1.350347e-07, -2.643895e-08, -5.110513e-08, 2.402032e-09, 7.433475e-08, 
    -3.047597e-08, -5.280697e-09, 5.616536e-08, -1.206477e-08, -9.795997e-09, 
    5.17332e-09, -8.847816e-08, 3.727081e-08, -6.911307e-09, -8.934251e-09, 
    1.870902e-07, 3.093828e-07, 3.661449e-08, -1.564176e-07, 2.455369e-08, 
    -2.430664e-08, -1.390248e-07, 4.746425e-11, -1.484085e-07, -2.422786e-08, 
    2.493009e-08, -2.157982e-08, 3.662916e-08, 4.702031e-09, -2.618168e-08, 
    1.121836e-07, -3.695875e-08, -1.065459e-10, -1.45414e-09, -3.038173e-08, 
    -3.772931e-08, -6.1202e-08, -2.792291e-08, 2.409928e-08, 1.799509e-08, 
    -2.373838e-09, -7.445067e-09, -2.134499e-08, -5.403598e-08, 
    -1.536762e-09, -1.431931e-09, 1.24937e-08, -1.31644e-09, -4.235829e-10, 
    -7.822285e-08,
  1.203773e-08, -1.973945e-09, -7.840299e-09, -4.070898e-09, 1.16089e-08, 
    2.87821e-08, 6.797575e-08, 7.12123e-09, -4.399931e-08, -4.261665e-09, 
    3.29419e-09, -6.755272e-10, -4.327683e-08, -1.500064e-08, 1.115507e-08, 
    -4.745196e-09, -6.134739e-08, 6.08037e-09, -2.022965e-08, -5.834863e-09, 
    1.559442e-09, 6.977314e-08, -9.122232e-10, 1.007038e-09, -3.781543e-08, 
    -2.640795e-07, 2.085108e-08, 2.13638e-08, -6.2141e-08, -1.650703e-07, 
    2.930244e-08, -7.948813e-08, 1.641536e-08, 5.826007e-08, -1.322933e-07, 
    2.486058e-08, 9.900385e-09, 2.143432e-08, 1.110449e-07, 2.447183e-07, 
    1.110886e-07, 3.270657e-09, 2.234052e-08, -3.710695e-08, 3.280365e-08, 
    -1.516295e-07, 2.087136e-07, 2.698314e-07, -8.343515e-08, -1.1e-08, 
    -1.670327e-08, -4.988112e-08, -5.082005e-08, 2.82987e-09, 4.210737e-08, 
    -1.000444e-09, 5.245397e-08, 1.914187e-08, 9.382367e-08, 3.272973e-08, 
    2.514867e-09, 5.308721e-09, 1.747242e-08, -2.983138e-08, -4.682772e-08, 
    2.666172e-08, 7.323274e-08, 3.415869e-08, 1.81343e-08, 2.564911e-08, 
    2.411044e-07, -5.288848e-08, -8.511347e-08, -8.868369e-09, 7.344475e-08, 
    -2.190188e-08, -8.456539e-09, 3.878077e-08, -1.171774e-08, -1.700982e-08, 
    2.820002e-09, -5.341139e-08, 5.880491e-08, -2.224813e-07, -2.616468e-08, 
    2.289592e-07, 1.908554e-07, 6.153493e-08, -1.792387e-07, 2.779041e-08, 
    3.946184e-09, -1.678654e-07, -7.890151e-10, -1.450485e-07, -3.5433e-08, 
    8.57847e-08, -9.470341e-09, 3.897833e-08, 4.157187e-09, -2.371289e-08, 
    4.28216e-07, -2.922133e-08, -4.081706e-09, 3.368683e-11, 3.050218e-10, 
    -4.507081e-08, -3.308946e-08, -1.893818e-08, 3.668151e-08, 1.935871e-08, 
    -6.136361e-09, -5.927518e-09, -1.876992e-08, -5.416723e-08, 
    -1.936883e-09, -1.308558e-09, 1.228078e-08, -1.318224e-09, -6.214265e-10, 
    -9.215967e-08,
  -4.306116e-09, -5.593051e-09, 1.200908e-08, 2.317222e-08, 7.52982e-09, 
    2.897866e-08, 8.431959e-08, 4.617607e-08, -1.629667e-08, -1.704882e-08, 
    9.432938e-09, -9.319217e-08, -4.227979e-08, -5.653021e-08, 1.039905e-08, 
    -5.475663e-09, -3.839709e-08, 7.145752e-08, 5.126992e-10, -5.285494e-08, 
    2.358354e-08, -2.072045e-08, -5.870447e-09, 1.237936e-09, -4.385345e-08, 
    -1.567749e-07, 1.807973e-08, 1.508658e-08, -3.604544e-08, -1.972932e-07, 
    2.632339e-08, -1.149823e-07, 1.892317e-09, 2.51656e-08, -1.27072e-07, 
    5.114657e-09, -1.841113e-09, 2.058312e-08, 1.106999e-07, 2.770363e-07, 
    4.438086e-08, -4.494609e-09, 1.603161e-08, -3.793755e-08, 1.561614e-08, 
    -1.33571e-07, 1.550218e-07, 3.459192e-07, -7.627134e-08, -9.849032e-09, 
    -1.029699e-08, -3.947218e-08, -6.72657e-08, 1.019482e-08, 2.445582e-08, 
    -8.838015e-10, 4.301398e-08, 1.935885e-08, 1.267506e-07, -1.553946e-08, 
    3.053287e-09, -5.621928e-09, -6.716357e-08, -3.603547e-08, -2.916761e-08, 
    2.115701e-08, 6.254402e-08, 3.370008e-08, 2.589275e-08, 1.059163e-08, 
    3.820595e-07, -8.877089e-08, -4.328774e-08, -2.881848e-09, 6.568937e-08, 
    -6.637379e-09, -1.107e-08, 2.371814e-08, -5.78566e-09, -2.769673e-08, 
    -4.686171e-10, -6.669257e-09, 6.522669e-08, -1.62583e-07, 2.953777e-08, 
    1.230375e-07, -1.043621e-07, 9.402049e-08, -2.105703e-07, -1.485409e-08, 
    1.884121e-08, -1.512634e-07, -1.997023e-09, -1.805974e-07, -5.984259e-08, 
    9.698289e-08, 5.824593e-08, 1.396245e-08, 5.837819e-10, -2.084792e-08, 
    1.993272e-07, -1.204982e-08, -8.853078e-09, -3.180816e-10, -1.575074e-08, 
    -3.541197e-08, -2.40982e-09, 1.468777e-08, 3.569869e-08, 1.27601e-08, 
    -1.792375e-08, -3.924129e-09, 1.287049e-09, -5.23022e-08, -2.259753e-09, 
    -9.796167e-10, 7.55e-09, -1.228713e-09, -6.99373e-10, -1.517034e-07,
  -1.373257e-08, -1.445676e-08, 1.331659e-08, 2.669083e-08, 5.201855e-09, 
    2.27493e-08, 9.039491e-08, 6.185803e-08, 1.024841e-08, -2.728143e-09, 
    3.498144e-10, -1.479411e-07, -1.861281e-09, -7.076994e-08, 1.289345e-08, 
    -3.323848e-10, -3.47031e-08, 8.44052e-08, -2.499891e-08, -1.897251e-08, 
    1.741894e-07, 8.482323e-08, -1.541962e-07, -3.000105e-08, -2.507386e-08, 
    -8.217944e-08, 1.143837e-08, 1.346405e-08, -1.284616e-08, -2.301522e-07, 
    4.22998e-08, -1.173612e-07, -4.860567e-09, -4.699905e-08, -1.196945e-07, 
    -2.981665e-09, -1.825231e-08, 1.902404e-08, 1.082143e-07, 3.093996e-07, 
    -1.225842e-08, 1.528227e-07, -2.223639e-07, -2.537994e-08, 2.631168e-08, 
    -8.793813e-08, 3.123768e-07, 3.781767e-07, -5.826903e-08, -6.908628e-09, 
    -3.571074e-09, 2.267939e-09, -9.797213e-08, 9.467954e-09, 9.788221e-09, 
    -6.394373e-09, 4.74987e-08, -4.31503e-09, 1.251811e-07, -1.650066e-08, 
    -2.81716e-10, -5.723177e-08, -1.317221e-08, -5.461594e-08, 6.408003e-09, 
    2.563411e-09, 2.600211e-08, 4.111462e-08, 1.576541e-08, -7.312678e-09, 
    1.675365e-07, 4.982178e-08, -1.153091e-08, -5.378183e-09, 3.988346e-08, 
    -1.305898e-08, -4.516224e-09, 1.848869e-08, -1.662426e-09, 1.526167e-07, 
    -3.275375e-09, 3.938e-08, 5.811296e-08, -7.448602e-08, 9.638916e-08, 
    4.59014e-08, -2.792896e-07, 9.128712e-08, -2.497324e-07, -7.668172e-08, 
    -1.13755e-08, -1.180173e-07, -1.100119e-09, -2.170563e-07, -5.40814e-08, 
    4.295648e-08, 1.135358e-07, -2.261663e-08, -1.174965e-08, -3.473242e-08, 
    -6.226662e-08, -2.048949e-09, -8.544482e-09, -2.833843e-09, 
    -1.474996e-08, -1.690046e-08, 2.570471e-08, 4.928984e-08, 2.418039e-08, 
    8.319603e-10, -3.539446e-08, -4.94731e-09, 1.392584e-08, -3.094158e-08, 
    -2.394813e-09, -1.426349e-09, 1.012391e-08, -1.237616e-09, -7.761898e-10, 
    -1.759391e-07,
  -1.711862e-08, -2.813397e-08, -9.832888e-09, 3.139235e-09, 4.190383e-09, 
    1.423871e-08, 7.720234e-08, 5.034065e-08, 1.645765e-08, 9.140535e-09, 
    -5.456957e-08, -7.103847e-08, 3.674415e-08, -4.650303e-08, -6.172161e-08, 
    5.392238e-09, -4.156077e-08, 3.794241e-08, -3.907371e-08, -7.140386e-08, 
    1.393261e-07, 1.31285e-07, -9.976441e-08, 1.448882e-08, -5.536663e-09, 
    -6.586845e-08, -7.035055e-09, 1.500246e-08, -3.923674e-09, -2.296212e-07, 
    -9.317887e-09, -6.794414e-08, -6.761979e-09, -4.549963e-08, 
    -1.285811e-07, -8.599159e-09, -3.563277e-08, 1.823719e-08, 1.005461e-07, 
    3.316874e-07, -1.976816e-08, 3.534785e-08, -2.274628e-07, -1.36616e-08, 
    -1.618116e-08, -4.388232e-08, 3.222244e-07, 3.365508e-07, -4.02282e-08, 
    -6.1452e-09, 1.806285e-09, 5.67411e-10, -1.662276e-07, 1.155152e-08, 
    -3.168884e-09, -1.059459e-08, 4.965784e-08, -2.525687e-08, 7.728204e-08, 
    5.164443e-08, -4.885919e-09, -1.092227e-07, 3.735352e-08, -1.459705e-08, 
    2.401573e-08, -2.439299e-08, 8.933398e-09, 3.656839e-08, 2.032868e-08, 
    -1.280171e-08, 1.398806e-07, 1.59008e-07, -2.632476e-08, -2.430363e-08, 
    1.202598e-08, -1.918238e-09, 4.379788e-08, 1.19179e-08, -4.330491e-09, 
    -1.116439e-08, 1.398121e-09, 4.648207e-08, 3.764706e-08, -6.236212e-08, 
    1.410389e-07, -5.25082e-08, -2.283199e-07, 2.792524e-08, -2.584189e-07, 
    -7.217227e-08, -7.976371e-08, -1.0646e-07, 4.193964e-09, -2.607532e-07, 
    -7.28495e-08, 5.507375e-08, 5.372911e-08, 1.136357e-08, -2.659851e-08, 
    -6.344023e-08, -9.925486e-08, 5.69085e-09, -7.614744e-09, -5.903956e-09, 
    -5.154448e-09, -3.61398e-08, 1.019691e-08, 3.769162e-08, 9.220798e-09, 
    -1.132764e-08, -4.248011e-08, -2.443915e-08, 8.587563e-09, 1.418027e-08, 
    1.887577e-08, -8.609049e-10, 1.035394e-08, -1.2218e-09, -7.299406e-10, 
    -9.867688e-08,
  -2.56739e-09, -4.807544e-08, -6.780999e-08, -1.328544e-08, 1.731587e-08, 
    1.07168e-08, 5.564493e-08, 1.546778e-08, 1.226954e-08, 7.266181e-09, 
    -9.615371e-08, 3.261516e-08, 4.382059e-08, -4.836465e-09, -1.668434e-07, 
    5.08409e-09, -3.675342e-08, 2.301681e-08, -4.463318e-08, -7.572817e-08, 
    2.223544e-08, 9.264375e-08, -2.530226e-08, 8.806046e-08, 7.510721e-09, 
    -4.373032e-08, -8.686811e-10, 1.673732e-08, 1.291255e-09, -2.183228e-07, 
    -1.366857e-09, -3.234049e-08, 8.212396e-09, -1.075296e-08, -1.159765e-07, 
    -1.623721e-08, -4.925596e-08, 1.975025e-08, 9.281086e-08, 3.250722e-07, 
    2.628158e-08, -2.142417e-08, -7.291976e-08, -1.835287e-09, -2.605634e-08, 
    -1.345381e-08, 2.81971e-07, 2.505738e-07, -2.742149e-08, -1.360625e-09, 
    5.74164e-09, -2.569459e-07, -2.477579e-07, 1.603919e-08, -1.719809e-08, 
    -5.331856e-09, 3.360299e-08, -4.473031e-08, 4.805447e-08, -1.47716e-08, 
    -6.622599e-09, -1.124653e-07, 1.106024e-07, 2.997831e-08, 1.684321e-08, 
    -4.045364e-08, 3.330581e-08, 3.31396e-08, 1.302863e-08, 1.718945e-08, 
    1.17313e-07, 1.68353e-07, -6.640369e-08, -6.284756e-08, -6.93492e-08, 
    7.124072e-09, 3.706158e-08, 1.58698e-08, 2.396299e-09, -7.743483e-08, 
    -7.204903e-09, 4.822623e-08, 1.342005e-08, -6.899188e-08, 2.386673e-07, 
    -7.37316e-08, -9.06233e-08, -1.133822e-08, -2.246208e-07, 3.390198e-09, 
    -3.012888e-07, -1.097715e-07, 1.324395e-09, -2.991605e-07, -2.2378e-08, 
    6.097391e-08, -6.780685e-08, -1.702347e-09, -1.376293e-08, -4.732044e-08, 
    -2.901459e-08, -2.211066e-08, -6.210882e-09, -7.194295e-09, 4.246192e-08, 
    -8.140478e-08, -5.40424e-08, 2.089337e-09, -3.705964e-09, -1.965498e-08, 
    -3.532318e-08, -1.066983e-07, -4.075821e-08, 8.310394e-09, 8.111363e-08, 
    -1.877879e-10, 9.151307e-09, -1.873193e-09, -6.066116e-10, 3.784862e-08,
  -1.026509e-07, -8.426758e-08, -9.91393e-08, -1.661675e-08, 3.380632e-08, 
    1.518828e-08, -4.946031e-08, -6.95623e-08, -1.609561e-08, -6.309398e-08, 
    -8.580236e-08, -4.370673e-08, -6.198945e-09, -1.836662e-08, 
    -2.216894e-07, 2.690266e-08, -3.392221e-08, 1.18028e-08, 4.516646e-08, 
    -6.815543e-08, -5.624594e-08, 4.096279e-08, 9.204615e-08, 8.126e-08, 
    -7.188947e-08, 1.537245e-08, 5.859135e-09, 1.895779e-08, 5.763354e-10, 
    -2.080147e-07, 9.324879e-09, -2.798737e-08, 1.711675e-08, 8.708582e-09, 
    -1.497762e-08, -2.048495e-08, -5.537887e-08, 2.425728e-08, 1.454965e-07, 
    2.914413e-07, 4.870309e-08, -3.467159e-08, -1.175906e-08, 1.41334e-08, 
    -3.499969e-08, -1.84138e-08, 1.70797e-07, 1.860599e-07, -2.471262e-08, 
    2.462791e-09, 8.494339e-09, -1.566866e-07, -2.976516e-07, 1.939708e-08, 
    -2.609541e-08, -1.847241e-09, 1.704922e-08, -5.807114e-08, 7.528892e-08, 
    -6.738267e-08, -9.728751e-10, 1.00128e-08, 1.076293e-07, 6.248113e-08, 
    -1.381535e-08, -3.992017e-08, 5.782914e-08, 7.208433e-08, 8.339669e-09, 
    3.55771e-08, 8.292437e-08, 8.392198e-08, -7.138857e-08, -6.957106e-08, 
    6.504017e-09, 3.994688e-08, -1.18583e-08, 9.314277e-09, 5.270332e-09, 
    -4.081443e-08, -6.861569e-10, 5.435948e-08, -1.047511e-08, -7.66351e-08, 
    5.596468e-08, -8.398803e-08, -2.705741e-08, -1.501343e-08, -1.668893e-07, 
    6.966582e-08, -2.833448e-07, -1.115332e-07, 8.782877e-10, -2.874052e-07, 
    1.018719e-08, 4.859931e-08, -1.520982e-07, -8.268955e-09, 8.451877e-09, 
    -1.798072e-08, -4.89967e-08, 5.395509e-08, -5.305253e-09, -5.903836e-09, 
    6.541023e-08, -8.780495e-08, -9.684942e-08, -1.989309e-08, -1.98084e-08, 
    -2.363134e-08, -2.695316e-08, -4.327813e-08, -1.238909e-07, 1.114643e-09, 
    5.438307e-08, -1.782837e-10, 7.573774e-09, -2.021679e-09, -5.187957e-10, 
    3.929046e-08,
  -4.583632e-07, -1.391349e-07, -7.827572e-08, -7.095935e-09, 2.974087e-08, 
    9.411059e-08, -2.46158e-07, -2.183808e-07, -5.874057e-08, -5.631949e-08, 
    1.935803e-09, -2.916187e-08, -1.059112e-08, -1.322125e-07, -1.787486e-07, 
    5.224982e-08, -3.872547e-08, 2.042384e-08, 1.729069e-08, -1.695156e-08, 
    -5.07485e-08, 3.166804e-09, 7.83462e-08, 1.041138e-08, 6.888723e-08, 
    8.116086e-08, -2.621601e-08, 1.015388e-08, 2.81517e-09, -1.905747e-07, 
    5.962949e-08, -3.389306e-08, -1.30953e-08, 9.645021e-09, -1.656718e-08, 
    -2.211544e-08, -5.348963e-08, 2.724883e-08, 3.735981e-07, 2.401821e-07, 
    4.699672e-08, -1.649191e-07, 7.42638e-08, 3.223496e-08, 1.569782e-08, 
    -3.246436e-08, 8.080804e-08, 1.230467e-07, -2.287244e-08, 3.927212e-09, 
    1.03656e-08, -6.857266e-08, -2.747748e-07, 1.83975e-08, -3.449293e-08, 
    -1.930005e-09, 1.45813e-08, -1.470013e-08, -5.303596e-08, -4.833595e-08, 
    -7.598493e-08, 4.542079e-08, 4.570154e-09, 6.878406e-08, -4.042996e-08, 
    -3.973656e-08, 6.69167e-08, 1.010401e-07, -4.504898e-09, 4.816906e-08, 
    5.246335e-08, -4.542034e-08, -7.422858e-08, -7.730949e-08, 6.062704e-08, 
    5.341673e-08, -4.858927e-08, 8.834661e-09, -4.18612e-09, 9.814016e-10, 
    1.049648e-08, 6.853589e-08, -1.126983e-08, -1.043633e-07, -4.070688e-08, 
    -9.378203e-08, -2.517885e-08, -9.576581e-09, -6.038569e-08, 1.108584e-07, 
    6.721342e-08, -1.062279e-07, 7.18083e-09, -2.318562e-07, 4.970212e-08, 
    7.915167e-08, -1.192533e-07, 1.115581e-08, 1.722827e-08, -3.128854e-08, 
    -6.872136e-08, 4.386738e-08, -5.414677e-09, -4.45737e-09, 5.741816e-08, 
    -4.737961e-08, -1.358341e-07, -3.82376e-08, -3.284077e-08, -2.972143e-08, 
    -2.198095e-08, -3.67271e-09, -3.405427e-08, 2.169543e-09, 2.072073e-08, 
    -4.144113e-10, 6.302571e-09, -2.445407e-09, -4.089742e-10, -3.643385e-08,
  1.10898e-07, -1.811076e-07, -5.018012e-08, 1.503054e-09, 8.848394e-08, 
    7.459482e-08, -1.917425e-07, -1.576258e-07, -9.587995e-08, -1.506316e-08, 
    3.044585e-07, 1.033925e-08, 5.332936e-09, 8.896393e-08, -1.107461e-07, 
    7.605868e-08, -4.832944e-08, 4.064736e-08, 8.842449e-09, -2.819081e-08, 
    -3.851767e-08, 1.38765e-08, -2.717081e-08, -1.405748e-07, 8.975428e-08, 
    1.337943e-07, -7.076744e-08, 2.001229e-09, 1.230944e-08, -1.667498e-07, 
    5.929121e-08, -3.271805e-08, -3.267394e-08, 1.77746e-08, 3.914363e-08, 
    -4.210699e-08, -3.955756e-08, 2.712912e-08, 3.203778e-07, 1.8579e-07, 
    6.73768e-08, -1.99388e-07, 1.197011e-07, 4.817973e-08, 1.505498e-08, 
    -5.453114e-08, -6.615062e-08, 5.443746e-08, -7.037511e-09, 4.156306e-09, 
    1.183409e-08, -4.894707e-08, -2.6963e-07, 1.735486e-08, -4.33295e-08, 
    -9.803216e-10, 2.245167e-08, 1.639494e-07, -3.500749e-08, -4.393385e-08, 
    5.768482e-08, 1.300215e-07, -1.196319e-07, 6.511547e-08, -5.934391e-08, 
    -3.669663e-08, 7.0699e-08, 9.078701e-08, -1.317937e-08, 1.126162e-07, 
    2.710692e-08, -6.090534e-08, -1.071877e-07, -6.091989e-08, 5.774768e-08, 
    4.092283e-08, -4.401949e-08, 1.395546e-08, -7.952207e-09, -1.112084e-07, 
    1.060062e-08, 6.707135e-08, 1.513854e-09, -5.619188e-08, -1.326529e-07, 
    -9.477651e-08, -4.957667e-08, 9.54401e-10, 5.38285e-08, 1.145916e-07, 
    1.342494e-08, -1.13081e-07, 2.843649e-09, -1.368451e-07, 1.500597e-07, 
    2.134172e-07, -8.489112e-08, 1.257403e-07, 1.661567e-08, -3.582272e-10, 
    -5.728646e-08, 3.54883e-08, 4.614962e-08, -3.00804e-09, -4.903313e-10, 
    -2.296167e-08, -1.476839e-07, -7.095639e-08, -5.167965e-08, 
    -4.017954e-08, -2.117565e-08, -4.086246e-09, 1.461672e-09, 2.231786e-09, 
    -3.954369e-09, -5.801212e-10, 6.206619e-09, -2.557854e-09, -3.51065e-10, 
    -4.980586e-08,
  1.567047e-07, -1.982903e-07, -1.459583e-07, 2.113717e-08, 1.295799e-07, 
    1.770155e-08, -6.462182e-08, -5.489591e-08, -3.746908e-08, 1.69919e-07, 
    2.334505e-07, 2.620574e-07, 2.118446e-08, 1.237136e-07, 1.014964e-07, 
    9.321559e-08, -1.198809e-07, 4.018494e-08, 2.194429e-08, -6.029933e-08, 
    -7.831488e-09, 4.035104e-08, -5.149485e-08, 8.401855e-09, 1.495053e-07, 
    -9.399912e-09, -6.669273e-08, 2.173311e-08, 1.949076e-08, -1.443551e-07, 
    4.323175e-08, -4.883049e-08, -2.327891e-08, -9.010307e-09, 7.131547e-08, 
    -2.733219e-08, 5.859973e-08, 2.600046e-08, 2.647139e-07, 1.142152e-07, 
    9.644076e-08, -9.336662e-08, 1.466813e-07, 6.78672e-08, -1.765278e-08, 
    -7.857847e-08, -1.415676e-07, -1.079604e-08, -6.213815e-09, 3.847433e-09, 
    1.302494e-08, -1.077628e-07, -2.569382e-07, 2.180415e-08, -4.155588e-08, 
    -1.241062e-09, 1.880716e-08, 1.918508e-07, -1.851402e-08, -3.567239e-08, 
    1.274401e-08, 6.025897e-08, 3.906138e-08, 7.257669e-08, -8.080334e-08, 
    -2.265602e-08, 3.354336e-08, 2.685073e-08, -1.867335e-08, 6.016143e-08, 
    1.714358e-08, 3.508745e-08, -6.684189e-08, 2.919404e-08, 3.094809e-08, 
    2.365022e-08, -2.822196e-08, 4.895639e-09, -1.674078e-08, -9.608954e-08, 
    1.868671e-08, 7.469086e-08, 6.008082e-08, -7.210173e-08, -1.165697e-07, 
    -5.070973e-08, -5.230373e-08, 1.046391e-08, 1.351434e-07, 9.963952e-08, 
    -4.031205e-08, -1.086485e-07, 2.653877e-09, -5.103709e-08, 1.009051e-07, 
    6.323117e-08, -2.751776e-09, 1.156212e-07, 9.960502e-09, 8.302688e-08, 
    -4.379848e-08, -2.085599e-09, 1.490354e-07, -2.040323e-10, 3.00119e-08, 
    1.224606e-08, -1.50764e-07, -1.040027e-07, -7.391458e-08, -3.620931e-08, 
    -2.186147e-08, -1.980027e-09, 1.929209e-09, 2.570744e-09, -7.59934e-09, 
    -6.749474e-10, 8.341033e-09, -2.41031e-09, -4.880718e-10, -2.987821e-08,
  2.231248e-07, -1.900831e-07, -4.970086e-07, 1.765051e-08, 5.183807e-08, 
    -4.302086e-08, -3.327233e-08, -1.268324e-07, 5.427802e-08, 7.204216e-08, 
    -1.147038e-08, 2.551328e-07, 1.578346e-07, 8.399633e-08, 5.419412e-08, 
    1.099926e-07, -1.071988e-07, 4.183414e-08, -2.000746e-10, -9.082709e-08, 
    -1.804193e-08, 1.412962e-07, -4.330167e-08, -2.99197e-08, 1.0871e-07, 
    -2.588155e-08, -4.813779e-08, 2.618077e-08, 2.497967e-08, -1.731933e-07, 
    8.301873e-08, -5.565897e-08, 1.727545e-08, -2.50763e-08, -5.204669e-08, 
    -3.704855e-08, 1.551901e-07, 2.34687e-08, 1.97264e-07, 2.613569e-08, 
    1.118695e-07, -1.549432e-07, 5.886818e-08, 6.390257e-08, -3.27687e-08, 
    -7.996738e-08, -1.36995e-07, -5.096314e-08, -1.399438e-08, 2.532914e-09, 
    1.369092e-08, -2.255696e-07, -1.271946e-07, 1.937789e-08, -4.34277e-08, 
    1.317403e-09, 3.269821e-08, -1.9114e-08, -2.168687e-08, -3.357317e-08, 
    1.345751e-08, 1.9673e-08, 4.309885e-08, 9.848353e-08, -6.026104e-08, 
    1.179245e-08, -8.517986e-10, -1.571203e-08, -1.647703e-08, 2.15295e-08, 
    1.865232e-08, 3.756696e-08, -7.849809e-08, -6.471208e-08, 1.637184e-08, 
    1.510733e-08, -8.752465e-09, 1.412707e-08, -3.611586e-08, -4.964312e-08, 
    2.096829e-08, 8.274726e-08, 4.429097e-08, -1.220672e-07, -3.209362e-08, 
    -1.48795e-08, 6.293425e-08, 8.296126e-09, 1.684413e-07, 7.801526e-08, 
    -9.327385e-08, -9.108368e-08, -2.258332e-09, 1.969403e-08, 8.769979e-08, 
    2.20478e-08, 2.292075e-09, 6.509225e-08, 1.222253e-08, 7.968161e-08, 
    -2.170913e-08, -2.825618e-08, 7.128209e-08, 4.404647e-09, 3.498229e-08, 
    1.077291e-08, -1.582993e-07, -1.225275e-07, -7.462057e-08, -2.673306e-08, 
    -2.224414e-08, -1.303931e-09, 4.094261e-09, 3.143043e-09, -7.963592e-09, 
    -8.951247e-10, 1.055059e-08, -2.349267e-09, -4.154685e-10, 1.035203e-07,
  2.230763e-07, -2.722443e-07, -5.030491e-07, -3.337755e-08, 1.031386e-07, 
    1.423587e-09, -1.730086e-08, 3.54554e-08, 3.82496e-08, 6.983157e-08, 
    -3.941307e-08, 2.510524e-07, 1.137428e-07, -1.281001e-08, -1.972614e-08, 
    1.147073e-07, -2.033093e-07, 4.260875e-08, -2.839434e-08, 1.855576e-07, 
    -3.828075e-08, -1.796377e-08, -1.701369e-08, -4.413005e-08, 5.43539e-08, 
    -3.652224e-08, 7.140659e-08, 2.378351e-08, 4.561093e-08, -1.656368e-07, 
    1.990463e-08, -2.600359e-08, 3.695402e-08, -1.009133e-07, 3.285561e-08, 
    -2.930938e-08, 1.976858e-08, 1.933178e-08, 6.649805e-08, -2.332705e-08, 
    1.498258e-07, -6.620803e-08, 5.238292e-09, 5.85082e-08, -4.405274e-08, 
    -8.10054e-08, -1.110345e-07, -5.295502e-08, -1.357848e-08, 8.813146e-10, 
    1.418975e-08, 2.598756e-08, -8.673769e-08, 2.419968e-08, -3.763192e-08, 
    9.69294e-10, -3.422224e-08, -2.938007e-08, -2.287748e-08, -4.990848e-08, 
    4.328808e-08, 2.400873e-08, 7.769711e-08, 1.055197e-07, -1.604653e-08, 
    2.074887e-08, -4.956291e-09, -6.394498e-08, -1.679371e-08, 1.683532e-08, 
    7.944664e-08, 1.132162e-08, 1.623354e-07, -5.042739e-08, 7.239009e-09, 
    -3.490186e-10, 3.111182e-08, -1.564501e-08, -1.859831e-08, -9.549717e-08, 
    2.001644e-08, 9.229628e-08, 2.786152e-08, 1.014763e-07, -4.008496e-08, 
    -6.338871e-08, 2.4145e-07, -3.733589e-08, 1.798853e-07, 6.123901e-08, 
    5.202196e-09, -6.83324e-08, -1.442095e-08, 1.000557e-07, 4.983258e-08, 
    1.308031e-09, -1.52741e-08, 2.184868e-08, 8.126335e-09, -2.263005e-08, 
    3.368768e-09, 2.474481e-08, 3.995981e-08, 7.090726e-09, 2.332001e-08, 
    -2.620936e-08, -1.604906e-07, -1.329593e-07, -7.181768e-08, 
    -2.091474e-08, -2.123397e-08, 6.028813e-10, 6.20139e-09, 3.680952e-09, 
    -8.263328e-09, 4.044864e-10, 3.462247e-09, -2.087262e-09, -3.858602e-10, 
    -3.152297e-08,
  2.261561e-07, -6.654818e-08, 1.716705e-08, -2.022614e-08, 3.301614e-08, 
    4.259607e-08, 5.630341e-08, 4.89573e-08, 6.36453e-09, 2.482011e-09, 
    -8.445033e-08, 8.536631e-08, 9.616656e-09, -2.010552e-08, -2.763272e-08, 
    1.206832e-07, -1.222225e-07, 2.55294e-08, -1.004344e-07, -4.43697e-08, 
    -2.400589e-08, -4.351159e-08, -5.285187e-09, -5.064487e-08, 1.621095e-08, 
    -3.84548e-08, 1.07724e-07, 1.534102e-08, 1.18412e-07, -6.677828e-08, 
    6.627204e-08, 1.499416e-09, -8.49318e-08, -1.038277e-07, 5.175048e-08, 
    -1.839851e-08, -3.261326e-08, 1.520081e-08, -5.098491e-08, -4.161408e-08, 
    2.16156e-07, 4.714821e-09, -2.070226e-08, 2.841143e-08, -5.421691e-08, 
    -1.03667e-07, -6.086725e-08, -4.436583e-08, -2.202824e-08, 1.10343e-09, 
    1.467238e-08, 4.636149e-08, -6.918558e-08, 2.543641e-08, -2.238011e-08, 
    9.564474e-10, -1.340336e-07, -1.008278e-07, -2.259136e-08, -7.927461e-08, 
    6.314588e-08, 2.568061e-08, 7.737208e-08, 9.677369e-08, -9.927953e-08, 
    4.088042e-08, 2.069066e-08, -1.146969e-07, 2.456579e-08, -1.39039e-10, 
    4.818662e-08, -4.689844e-08, 2.37078e-08, -1.546971e-08, 2.60852e-09, 
    -1.647538e-08, -1.298037e-08, 8.279812e-10, -1.631051e-08, -4.512128e-08, 
    3.140394e-08, 9.438787e-08, 2.765108e-08, -2.936292e-08, -3.504374e-08, 
    -1.310269e-07, 3.330798e-07, -1.313169e-07, 1.940184e-07, 4.963783e-08, 
    2.530055e-08, -4.618396e-08, -8.330289e-09, 1.261439e-07, 3.049763e-09, 
    -5.919279e-09, -2.600893e-08, -2.07707e-08, 7.39476e-09, -2.918121e-08, 
    -2.482693e-09, -1.760099e-08, 5.511815e-09, 8.39519e-09, 4.748244e-09, 
    -6.10097e-08, -1.722849e-07, -1.383589e-07, -7.244773e-08, -1.977469e-08, 
    -2.459831e-08, 1.811827e-09, 7.267658e-09, 3.998366e-09, -9.097562e-09, 
    3.842615e-09, 5.813803e-09, -2.665157e-09, -5.169198e-10, -2.495176e-08,
  2.270633e-07, -2.799425e-08, 8.542429e-10, 1.74623e-09, 7.476046e-09, 
    2.374441e-08, 1.917442e-08, 2.546403e-08, -2.83012e-09, -1.135436e-08, 
    -2.489719e-08, -5.723268e-08, 1.119588e-09, -2.301749e-08, -2.956017e-08, 
    1.306694e-07, -9.958001e-08, 1.790261e-08, -1.912801e-07, -6.163418e-08, 
    -2.318416e-08, -5.743709e-08, 3.185278e-09, -5.345782e-08, -3.330797e-09, 
    -3.879904e-08, 4.498997e-08, 2.548813e-08, 1.700564e-07, -1.580747e-08, 
    2.041268e-07, -8.687266e-09, -9.728228e-08, -1.190492e-07, 1.883973e-08, 
    6.738674e-09, -3.851699e-08, 1.243063e-08, -2.176191e-07, -4.805845e-08, 
    2.48111e-07, 6.232767e-08, -3.059779e-08, 1.671303e-08, -8.236611e-08, 
    -1.170413e-07, -2.786089e-08, -3.658499e-08, -1.531312e-08, 3.416332e-09, 
    1.525524e-08, 5.707534e-09, -6.62594e-08, 2.869433e-08, -7.415464e-09, 
    1.901981e-10, -1.713433e-07, -1.635352e-07, -2.241646e-08, -3.772533e-08, 
    6.736514e-08, 2.427919e-08, 9.103337e-08, 9.520722e-08, -1.040386e-07, 
    9.183623e-10, 6.733831e-08, -1.877643e-07, 6.944288e-08, -3.494438e-08, 
    9.886207e-09, -1.660615e-07, -4.277013e-08, 1.70412e-08, -7.256169e-10, 
    -1.983904e-08, -1.49428e-08, 6.760843e-09, -9.806802e-09, -8.055054e-08, 
    1.717603e-08, 9.546776e-08, 2.742411e-08, -2.09659e-08, 3.523769e-08, 
    -1.332912e-07, 1.719939e-07, -1.378658e-08, 2.032514e-07, 4.235153e-08, 
    3.029868e-08, -5.400761e-08, -7.618723e-09, 1.317993e-07, -2.593652e-09, 
    -8.505232e-09, -5.211136e-08, -7.613153e-08, 1.891522e-08, 3.057993e-09, 
    -4.034132e-08, -1.729543e-08, -9.247984e-09, 8.697526e-09, -2.482193e-08, 
    -8.687334e-08, -2.086504e-07, -1.406777e-07, -7.314202e-08, 
    -1.986177e-08, -2.309366e-08, 1.275339e-09, 7.84371e-09, 4.655476e-09, 
    -7.544713e-09, 7.816698e-09, 1.998188e-09, -1.909058e-09, -6.07713e-10, 
    -2.341562e-08,
  2.237981e-07, -2.432512e-08, 3.186403e-08, 7.619178e-09, 7.565745e-09, 
    3.451044e-08, 2.150409e-08, 3.508262e-08, -8.082225e-09, -1.074807e-08, 
    -1.109743e-08, -7.409494e-08, -2.525326e-09, -2.328125e-08, 
    -3.017146e-08, 1.716907e-07, -5.598832e-08, 1.699794e-08, -1.296468e-07, 
    -6.471362e-08, -2.273384e-08, -6.316168e-08, 3.720743e-09, -5.598463e-08, 
    -1.003139e-08, -3.832656e-08, 1.653746e-08, 1.270671e-07, 5.138349e-08, 
    2.065675e-07, 8.95061e-08, 1.113333e-07, -1.472456e-07, -1.047052e-07, 
    1.047863e-08, 1.290607e-08, -4.055568e-08, 1.067758e-08, -2.312779e-07, 
    -5.168852e-08, 3.112865e-07, 8.586937e-08, -3.681922e-08, 1.500352e-08, 
    -9.215296e-08, -1.27187e-07, 5.849188e-11, -3.316649e-08, -1.595536e-08, 
    -2.517382e-10, 1.585025e-08, -4.412868e-09, -5.94337e-08, 3.365049e-08, 
    6.366079e-09, -1.679155e-10, -5.193056e-08, -1.770784e-07, -2.238705e-08, 
    -1.207e-08, 7.069298e-08, 2.243314e-08, 9.351299e-08, 8.803075e-08, 
    -8.85836e-08, -1.092776e-07, 3.735067e-09, -1.448681e-07, -2.416505e-08, 
    -1.391447e-08, 2.575928e-08, -1.966893e-07, -5.421782e-08, 1.752846e-08, 
    -3.217643e-09, -2.501508e-08, -1.524661e-08, 1.177679e-08, -7.404324e-09, 
    -1.433966e-08, -4.243299e-08, 1.0454e-07, 2.665593e-08, -2.170657e-08, 
    5.880304e-08, -7.753636e-08, 1.102086e-07, -3.232117e-10, 2.096701e-07, 
    3.856843e-08, 3.239552e-08, -6.803157e-08, -6.683507e-09, 1.229851e-07, 
    8.161896e-08, -1.037759e-08, -5.26908e-08, -3.763148e-09, 2.090144e-08, 
    -1.599706e-08, -5.376648e-08, -2.069243e-08, -5.738798e-08, 8.336528e-09, 
    2.362913e-08, -2.311765e-08, -2.561684e-07, -1.406721e-07, -7.275912e-08, 
    -2.068293e-08, -2.258048e-08, 1.998615e-10, 7.600647e-09, 5.285528e-09, 
    -3.450509e-09, 1.272983e-08, -7.754721e-10, -1.628777e-09, -5.20032e-10, 
    -2.20482e-08,
  2.287792e-07, -2.251528e-08, 6.045354e-09, 9.730741e-09, 8.455174e-09, 
    5.422231e-08, 2.082089e-08, 3.825193e-08, -1.02529e-08, -1.107475e-08, 
    -4.0896e-09, -7.948421e-08, -3.923503e-09, -2.383518e-08, -3.025144e-08, 
    2.116312e-07, -1.288845e-08, 1.042184e-08, -8.067285e-08, -6.590454e-08, 
    -2.255416e-08, -6.600868e-08, 2.08928e-09, -5.706039e-08, -1.505754e-08, 
    -3.833503e-08, 2.636847e-08, 1.693428e-08, 3.991937e-08, 4.485338e-08, 
    5.546968e-08, 7.463262e-08, 1.950508e-08, -6.259921e-08, 6.253856e-09, 
    1.401355e-08, -4.160736e-08, 8.827399e-09, -3.228511e-07, -5.319991e-08, 
    3.466078e-07, 1.013761e-07, -3.871642e-08, 1.889523e-08, 1.917664e-08, 
    -1.366748e-07, 7.132371e-09, -3.369834e-08, -1.579114e-08, -2.642409e-09, 
    1.640809e-08, -6.733728e-09, -5.441043e-08, 3.824986e-08, 1.137522e-08, 
    -1.435467e-09, -1.343534e-08, -1.861236e-07, -2.253522e-08, 5.478564e-08, 
    7.258785e-08, 2.179485e-08, 9.487832e-08, 8.671517e-08, -7.805353e-08, 
    1.241189e-07, -1.888401e-08, -1.281226e-07, -4.212865e-08, -4.701172e-08, 
    -2.139757e-09, -1.523838e-07, -6.645888e-08, 1.707753e-08, -4.796348e-09, 
    -3.635245e-08, -1.420183e-08, 1.433114e-08, -3.483454e-10, -2.407256e-08, 
    -2.223413e-08, 1.088744e-07, 2.636096e-08, -2.182054e-08, 7.100886e-08, 
    -8.240801e-08, 9.333411e-08, 2.354824e-08, 2.12246e-07, 3.814836e-08, 
    3.308315e-08, -6.186621e-08, -5.313524e-09, 1.122081e-07, 3.861697e-08, 
    -1.191561e-08, -5.431087e-08, -4.49449e-08, 2.123357e-08, -6.946277e-09, 
    3.403727e-09, -2.239241e-08, -7.805246e-08, 8.186674e-09, 1.101381e-08, 
    -3.040083e-08, -2.630792e-07, -1.33164e-07, -7.186139e-08, -2.22023e-08, 
    -2.262033e-08, 4.775416e-10, 7.984852e-09, 5.212371e-09, 3.987964e-09, 
    9.112114e-10, -3.240388e-09, -1.252555e-09, -4.689582e-10, -2.074097e-08,
  2.283649e-07, -2.056493e-08, 3.886839e-09, 1.156116e-08, 9.370069e-09, 
    6.015978e-08, 2.002355e-08, 3.948833e-08, -1.163903e-08, -1.135106e-08, 
    -1.202125e-09, -8.125517e-08, -4.265871e-09, -2.491674e-08, -3.00771e-08, 
    2.144398e-07, 2.110778e-09, 1.052678e-08, -5.521041e-08, -6.664777e-08, 
    -2.235242e-08, -6.617029e-08, -1.668354e-09, -5.715447e-08, -1.56997e-08, 
    -3.792309e-08, -1.065632e-08, 1.944682e-08, 3.84515e-08, 4.869764e-08, 
    4.666902e-08, 7.923791e-08, 8.728875e-10, -5.024231e-08, 4.370463e-09, 
    1.687374e-08, -4.225103e-08, 5.986536e-09, -3.210163e-07, -5.502585e-08, 
    4.284975e-07, 1.103791e-07, -3.955989e-08, 2.558123e-08, -8.91514e-08, 
    -1.306867e-07, 1.450775e-08, -3.53794e-08, -1.277081e-08, -2.196636e-09, 
    1.66368e-08, -7.635094e-09, -5.127371e-08, 3.862197e-08, 8.347055e-09, 
    -3.439766e-09, -3.459036e-09, -1.91304e-07, -2.293592e-08, 9.509742e-08, 
    7.322046e-08, 2.101524e-08, 9.203086e-08, 8.797981e-08, -4.894564e-08, 
    -6.148764e-08, -3.986304e-08, -1.027383e-07, -4.470371e-08, 
    -4.619051e-08, -3.72313e-09, -8.006759e-08, -6.898154e-08, 1.639376e-08, 
    -5.757226e-09, -5.329878e-08, -1.455662e-08, 1.635735e-08, 5.314453e-09, 
    -4.960384e-09, -8.02612e-09, 1.050013e-07, 2.610494e-08, -2.15623e-08, 
    7.936183e-08, -4.102969e-08, 8.197253e-08, 2.244394e-08, 2.132228e-07, 
    3.899657e-08, 3.255593e-08, -6.036803e-08, -3.197982e-09, 9.523244e-08, 
    4.140088e-08, -1.306816e-08, -5.4561e-08, -3.358241e-08, 2.04617e-08, 
    5.627953e-10, 2.004742e-08, -2.248508e-08, -9.085988e-08, 8.468341e-09, 
    1.084629e-08, -5.054471e-08, -2.258556e-07, -1.238237e-07, -7.136555e-08, 
    -2.464787e-08, -2.142724e-08, 2.192905e-09, 7.403514e-09, 5.893185e-09, 
    2.056561e-08, 2.946763e-10, -1.670912e-09, -9.653789e-10, -3.425598e-10, 
    -2.025706e-08,
  2.280213e-07, -1.893977e-08, -2.585921e-09, 1.492742e-08, 1.041985e-08, 
    6.367213e-08, 1.921853e-08, 3.939374e-08, -1.295609e-08, -1.126705e-08, 
    1.236913e-09, -8.117797e-08, -4.126264e-09, -2.511081e-08, -2.980357e-08, 
    1.596269e-07, 6.725838e-09, 1.101301e-08, -3.906635e-08, -6.708274e-08, 
    -2.213426e-08, -6.64329e-08, -5.235734e-09, -5.625736e-08, -1.628462e-08, 
    -3.707305e-08, -2.812283e-08, 9.175665e-10, 3.910714e-08, 6.06359e-08, 
    3.920741e-08, 3.818604e-08, -1.237083e-08, -6.460664e-08, 3.615469e-09, 
    7.483095e-09, -4.270861e-08, 2.601027e-09, -2.4824e-07, -5.528352e-08, 
    4.852027e-07, 1.139364e-07, -4.075378e-08, 1.732999e-08, -9.917233e-08, 
    -1.253686e-07, 1.71525e-08, -3.63074e-08, -1.069295e-08, -2.735007e-09, 
    1.705551e-08, -7.860308e-09, -4.939272e-08, 4.020901e-08, 6.565034e-09, 
    -2.198306e-09, -1.113938e-08, -1.940532e-07, -2.362939e-08, 8.325101e-08, 
    7.30771e-08, 1.997796e-08, 9.002383e-08, 8.829766e-08, -4.434846e-08, 
    -6.05753e-08, -1.280716e-08, -9.000189e-08, -1.104036e-08, -6.698076e-08, 
    -3.842058e-08, 5.770107e-08, -6.949904e-08, 1.538695e-08, -6.415373e-09, 
    -4.771857e-08, -1.430344e-08, 1.818063e-08, 1.06355e-08, -2.100251e-09, 
    -3.953176e-09, 9.975994e-08, 2.586989e-08, -2.075262e-08, 8.691791e-08, 
    -3.925072e-08, 7.788083e-08, 2.173317e-08, 2.076642e-07, 3.968438e-08, 
    3.224443e-08, -4.809995e-08, -8.376162e-10, 8.1458e-08, 3.041464e-08, 
    -1.397584e-08, -5.536535e-08, -4.976687e-08, 1.864646e-08, 4.695085e-09, 
    2.008687e-08, -2.239914e-08, -9.015213e-08, 8.27611e-09, 9.995688e-09, 
    -5.15663e-08, -1.763731e-07, -1.140589e-07, -7.106576e-08, -2.58608e-08, 
    -1.852288e-08, 3.085461e-09, 6.846676e-09, 6.978098e-09, 5.875063e-08, 
    -1.115973e-09, -3.373415e-09, -6.470557e-10, -4.283507e-10, -2.096021e-08,
  2.276668e-07, -1.669372e-08, -4.4883e-09, 1.671623e-08, 1.159816e-08, 
    6.634747e-08, 1.817801e-08, 3.966949e-08, -1.472739e-08, -1.255495e-08, 
    5.329696e-09, -7.837917e-08, -3.663843e-09, -2.34848e-08, -2.936082e-08, 
    1.054031e-07, 6.329366e-09, 1.00506e-08, -3.116331e-08, -6.721399e-08, 
    -2.219991e-08, -6.700333e-08, -5.717368e-09, -5.404257e-08, 
    -1.685311e-08, -3.625536e-08, -4.151678e-08, -1.525729e-08, 4.003965e-08, 
    6.657973e-08, 3.457245e-08, 1.868244e-08, -3.519227e-08, -9.988668e-08, 
    2.357581e-09, 9.382404e-09, -4.305509e-08, 1.695e-09, -1.216702e-07, 
    -5.515171e-08, 5.855397e-07, 1.144679e-07, -4.207493e-08, 1.614611e-08, 
    -9.621891e-08, -1.210827e-07, 1.759366e-08, -3.634923e-08, -1.225129e-08, 
    -2.896101e-09, 1.714987e-08, -7.930623e-09, -4.84057e-08, 4.576979e-08, 
    5.966953e-09, 2.081379e-09, -1.830546e-08, -1.944885e-07, -2.467934e-08, 
    7.147159e-08, 7.224463e-08, 1.829284e-08, 8.810508e-08, 9.402089e-08, 
    -4.45464e-08, -6.206488e-08, -1.197407e-09, -8.285809e-08, -9.781218e-09, 
    -7.611919e-08, -4.957457e-08, 6.086833e-08, -6.732347e-08, 1.411598e-08, 
    -7.009227e-09, -2.478993e-08, -1.397937e-08, 1.793074e-08, 1.260769e-08, 
    -2.953016e-10, -4.644676e-09, 9.437016e-08, 2.559585e-08, -1.943243e-08, 
    8.872036e-08, -3.798249e-08, 7.583088e-08, 2.138285e-08, 2.068118e-07, 
    3.981694e-08, 3.209169e-08, -4.192226e-08, 1.268063e-09, 6.828295e-08, 
    2.632174e-08, -1.477115e-08, -5.60277e-08, -6.016018e-08, 1.651648e-08, 
    4.118522e-09, 1.845882e-08, -2.228719e-08, -8.926318e-08, 8.129113e-09, 
    8.896166e-09, -5.342946e-08, -1.284812e-07, -1.109236e-07, -7.286798e-08, 
    -2.445114e-08, -1.429129e-08, 5.082654e-09, 6.130051e-09, 7.514757e-09, 
    1.166601e-07, -6.803476e-10, -5.408836e-09, -3.999148e-10, -3.147704e-10, 
    -2.120493e-08,
  2.273062e-07, -1.309121e-08, -3.294133e-09, 1.740392e-08, 9.534403e-09, 
    6.889758e-08, 1.67683e-08, 3.915312e-08, -1.569589e-08, -1.275754e-08, 
    7.828646e-09, -7.525142e-08, -2.560739e-09, -2.17662e-08, -2.855103e-08, 
    6.579268e-08, 5.846051e-09, 9.506778e-09, -2.849094e-08, -6.69566e-08, 
    -2.255348e-08, -6.749366e-08, -5.757954e-09, -5.192697e-08, 
    -1.696918e-08, -3.471627e-08, -4.530824e-08, -2.299629e-08, 4.06597e-08, 
    6.9024e-08, 3.511735e-08, 1.672021e-08, -4.9162e-08, -1.647743e-07, 
    6.368168e-10, 1.706672e-08, -4.334814e-08, 1.181391e-09, -4.31607e-08, 
    -5.442362e-08, 7.209092e-07, 1.120536e-07, -4.306858e-08, 1.462314e-08, 
    -8.906062e-08, -1.137578e-07, 1.602751e-08, -3.529749e-08, -1.346096e-08, 
    -6.930954e-09, 1.697484e-08, -7.986216e-09, -4.791089e-08, 4.589259e-08, 
    4.520197e-09, 2.34553e-09, -3.181805e-08, -1.943716e-07, -2.630034e-08, 
    5.861793e-08, 7.046327e-08, 1.554343e-08, 8.584067e-08, 1.001983e-07, 
    -3.591553e-08, -7.321336e-08, 7.251515e-10, -8.673811e-08, 1.044214e-10, 
    -8.666183e-08, -5.694955e-08, 5.888643e-08, -6.575323e-08, 1.251959e-08, 
    -7.798374e-09, -7.694496e-09, -1.375595e-08, 1.667908e-08, 1.947562e-08, 
    -3.231833e-09, -6.448374e-09, 8.925707e-08, 2.490435e-08, -1.782308e-08, 
    9.011973e-08, -3.924225e-08, 7.977025e-08, 2.076212e-08, 2.078833e-07, 
    4.016999e-08, 3.196652e-08, -3.717631e-08, 2.361389e-09, 5.820279e-08, 
    2.543158e-08, -1.554725e-08, -5.560716e-08, -6.449801e-08, 1.476775e-08, 
    4.452966e-09, 2.233384e-08, -2.204909e-08, -9.14094e-08, 7.987488e-09, 
    7.498272e-09, -5.439477e-08, 1.233589e-07, -1.173801e-07, -7.801367e-08, 
    -2.156145e-08, -9.772805e-09, 9.008829e-09, 5.52717e-09, 8.76986e-09, 
    1.597503e-07, -2.482147e-09, -5.311179e-09, -7.899459e-09, -1.091067e-09, 
    -2.109761e-08,
  2.267576e-07, -4.977778e-09, 8.669758e-10, 2.055594e-08, 1.328101e-08, 
    7.265282e-08, 1.39637e-08, 3.778757e-08, -1.658532e-08, -1.240551e-08, 
    8.474558e-09, -7.088443e-08, -2.490879e-10, -1.879528e-08, -2.657339e-08, 
    5.985378e-08, 5.709751e-09, 9.098017e-09, -2.193097e-08, -6.570997e-08, 
    -2.1711e-08, -6.628591e-08, -5.229936e-09, -4.988226e-08, -1.668548e-08, 
    -3.108971e-08, -5.000004e-08, -2.599575e-08, 4.052117e-08, 7.063068e-08, 
    2.413412e-08, 1.58376e-08, -5.725531e-08, -1.440441e-07, -2.215643e-09, 
    1.673754e-08, -4.362579e-08, 1.331884e-09, -8.263942e-08, -5.308391e-08, 
    9.785124e-07, 1.046645e-07, -4.430146e-08, 1.28287e-08, -7.901622e-08, 
    -9.996722e-08, 1.084368e-08, -3.277333e-08, -1.386245e-08, -6.907086e-09, 
    1.720355e-08, -8.159418e-09, -4.793882e-08, 4.642136e-08, 6.026795e-09, 
    1.100659e-09, -4.04367e-08, -1.761813e-07, -2.931759e-08, 4.816553e-08, 
    6.633945e-08, 1.043054e-08, 8.108952e-08, 1.099187e-07, -2.692002e-08, 
    -7.925917e-08, -9.473524e-10, -8.234429e-08, 4.463345e-09, -9.160806e-08, 
    -6.410437e-08, 5.853224e-08, -6.186019e-08, 9.490577e-09, -9.511474e-09, 
    -2.098682e-08, -1.275394e-08, 1.494323e-08, 1.971111e-08, 1.087756e-09, 
    -6.167113e-09, 8.263918e-08, 2.397695e-08, -1.48691e-08, 8.403458e-08, 
    -3.545574e-08, 7.136873e-08, 1.911212e-08, 2.090479e-07, 4.565209e-08, 
    3.031448e-08, -3.244168e-08, 3.314796e-09, 4.86735e-08, 2.5811e-08, 
    -1.641416e-08, -5.305242e-08, -5.960317e-08, 1.232047e-08, 5.536936e-09, 
    1.832143e-08, -2.12743e-08, -9.167398e-08, 7.780663e-09, 4.792241e-09, 
    -5.531115e-08, 1.756557e-07, -1.290307e-07, -8.455356e-08, -2.10955e-08, 
    -8.686129e-09, 1.008948e-08, 1.257763e-08, 1.056333e-08, 1.585975e-07, 
    -1.273554e-09, 9.760001e-09, 6.117713e-09, -2.600238e-09, -1.954641e-08,
  4.397412e-13, 5.126599e-13, 3.624884e-13, 1.103705e-13, -8.604897e-14, 
    -2.465141e-13, -1.693568e-13, 6.460755e-13, 4.084915e-13, 2.388562e-14, 
    -2.053231e-13, -4.3698e-13, -1.109027e-13, -1.620932e-13, -3.204268e-13, 
    5.236868e-13, -2.819949e-12, -8.03773e-13, -2.686899e-14, -5.277903e-13, 
    -4.036436e-12, -2.50922e-12, 4.300709e-13, -1.096233e-13, -1.058047e-12, 
    -1.284834e-13, 3.108537e-13, -7.418171e-14, 4.790371e-15, 3.562682e-15, 
    -1.259372e-13, 3.815215e-14, 1.043484e-13, 8.790787e-14, 3.433836e-13, 
    2.708602e-13, -1.153889e-12, 2.387904e-12, 3.246173e-13, 5.906273e-13, 
    7.883593e-13, 9.90815e-14, -1.898252e-14, -2.797476e-13, 1.690498e-13, 
    6.338985e-13, 1.882082e-12, 6.70305e-13, -7.748099e-13, 5.142734e-13, 
    2.985313e-13, 9.125167e-15, 3.642642e-12, -7.589868e-13, -5.402851e-14, 
    -8.546755e-13, 7.348956e-14, -3.37858e-13, 1.043058e-13, 2.414412e-12, 
    9.654479e-13, 5.751911e-14, 3.630173e-14, -3.103292e-12, -5.122798e-13, 
    -6.856759e-14, 3.468291e-13, -1.692108e-13, -2.076168e-13, -9.165292e-14, 
    2.780913e-13, 6.424071e-14, 1.740654e-13, 3.128125e-13, -3.896188e-13, 
    9.258653e-14, 4.703406e-13, -1.106299e-12, -1.80693e-12, -2.076451e-13, 
    8.647378e-14, 8.539541e-13, 2.408876e-13, -6.487749e-13, 6.831583e-13, 
    2.832302e-13, 1.364502e-13, -3.141006e-13, 8.373653e-13, 3.553701e-12, 
    1.869565e-14, 1.186176e-12, -4.170332e-13, 3.837538e-13, -1.412538e-13, 
    -3.286962e-13, 1.699092e-13, -6.550484e-13, 1.323381e-13, -4.184258e-13, 
    -1.173888e-12, 8.567684e-13, -1.203488e-12, -1.152974e-12, -6.286721e-14, 
    -1.088958e-13, -1.143209e-13, -1.275408e-12, -2.311395e-12, 
    -1.202055e-12, -6.078144e-13, -1.496194e-13, -6.537781e-14, -3.84863e-14, 
    6.266763e-13, -3.579057e-12, 2.832801e-12, -6.249623e-14, 1.87358e-13, 
    2.324984e-13,
  5.054852e-13, 4.126033e-13, 4.822647e-13, 5.546136e-13, 5.609583e-13, 
    5.022378e-13, 4.943824e-13, 4.394601e-14, 1.47295e-13, -1.601052e-13, 
    -1.189179e-13, 2.34393e-13, 3.69316e-14, -1.514697e-13, -3.081664e-13, 
    3.4179e-14, -2.337552e-13, 1.552181e-15, -4.404212e-14, -1.086153e-13, 
    -2.888105e-13, -8.117447e-13, -9.668546e-13, 2.317408e-14, -5.878176e-13, 
    -8.241824e-13, -8.765081e-13, -2.505759e-13, -2.609151e-13, 4.530134e-14, 
    1.651107e-13, -4.662652e-14, -1.102521e-14, -2.434069e-13, -2.449707e-13, 
    6.469594e-14, -3.522362e-13, 1.201316e-13, 1.678014e-13, 7.89599e-13, 
    -8.003102e-13, -6.245042e-14, -2.041199e-14, 1.159105e-13, -4.086312e-14, 
    9.146293e-14, -1.211118e-12, 1.560086e-13, -3.094822e-14, -3.622928e-14, 
    -7.098724e-14, -8.782405e-14, -6.201109e-13, 2.70903e-12, 1.054683e-13, 
    -1.759606e-12, 8.013738e-13, -1.664533e-12, -3.563461e-13, 1.653857e-12, 
    5.89028e-13, 2.031704e-13, -2.812191e-13, -2.147052e-13, -1.170473e-13, 
    9.935696e-14, 3.864834e-13, -7.295405e-14, -1.500417e-13, -3.363165e-13, 
    -1.237646e-12, 2.756771e-13, 1.664177e-13, -2.799327e-13, 1.638699e-12, 
    -1.570318e-12, -4.054329e-13, 1.37051e-12, -4.529126e-12, -8.892789e-13, 
    -2.088319e-13, -5.108691e-13, 1.72399e-12, -4.533228e-13, 7.392675e-13, 
    6.502777e-13, 5.072919e-13, 8.084023e-14, 9.674363e-13, -1.491746e-12, 
    1.981183e-13, -4.999747e-14, 7.479922e-14, 4.283975e-13, 1.940326e-13, 
    3.164216e-13, 2.48431e-13, 7.551587e-14, 2.63003e-13, 4.070509e-13, 
    -1.273604e-12, 5.602319e-13, 4.671504e-13, -3.932171e-12, -3.931278e-13, 
    1.836292e-13, 1.291191e-13, -1.318137e-13, 2.858137e-13, 5.907711e-13, 
    4.379027e-13, 5.312776e-13, 3.457767e-13, 1.468599e-13, 3.571627e-13, 
    9.037089e-14, -3.527348e-12, 1.47596e-12, -3.292708e-13, 4.604762e-13,
  -6.201983e-14, -1.607048e-14, -2.792211e-14, -1.21847e-13, -2.33577e-13, 
    -3.015505e-13, -2.041561e-13, 7.506495e-14, 1.933731e-13, 1.019462e-13, 
    2.350897e-14, -2.004091e-13, -3.830963e-13, -7.467638e-14, 1.049022e-13, 
    1.947331e-13, -1.661005e-13, -1.302916e-13, -4.275139e-13, -1.450604e-12, 
    -1.109141e-12, -1.638287e-12, -1.764505e-12, -5.272172e-13, 
    -9.452161e-13, -1.173783e-12, -3.484435e-13, -6.041001e-14, 
    -1.023764e-13, -5.170864e-14, 1.047357e-13, -1.249001e-16, -2.148282e-14, 
    -8.222589e-14, 4.911349e-14, 6.875056e-14, -7.996062e-13, -5.355091e-14, 
    1.366685e-13, -1.019956e-12, 7.514184e-13, 6.964568e-13, -6.40217e-14, 
    1.94636e-15, 4.971856e-13, 8.408552e-14, -1.865008e-12, -1.132528e-12, 
    1.564082e-13, 4.28082e-13, -5.821038e-14, -1.088879e-12, -4.088785e-13, 
    -2.815595e-11, 4.25493e-15, -9.670667e-13, -1.066772e-12, -1.651065e-12, 
    -1.911041e-12, 1.840765e-12, 3.889389e-13, -7.291945e-13, -8.830436e-14, 
    -1.210587e-13, -2.249562e-13, -2.570166e-14, -1.369599e-13, 
    -3.241851e-14, 1.321165e-13, -1.290495e-13, -4.543588e-14, 3.596567e-13, 
    5.398876e-13, -3.572698e-13, 3.73461e-13, -3.343811e-12, -5.883957e-13, 
    1.853968e-13, 2.397768e-12, -6.856044e-13, 9.891879e-13, 1.379515e-12, 
    -8.450463e-13, -4.520134e-13, -1.514899e-13, -6.319945e-13, 
    -1.970049e-12, 1.474515e-13, -1.388167e-12, -2.306932e-12, -2.397665e-13, 
    -1.426664e-13, 4.224607e-13, -3.573516e-12, -9.074685e-14, 9.246395e-13, 
    6.779966e-13, -7.69107e-14, 4.764938e-13, 2.966782e-12, 9.232753e-13, 
    -1.675075e-13, 6.019152e-13, -4.581752e-13, 4.967693e-13, 9.599127e-13, 
    1.035547e-12, 1.454489e-12, 1.176642e-12, 5.701412e-13, 6.013801e-13, 
    6.733364e-13, 8.444079e-13, 8.007345e-13, 5.88668e-13, 1.35981e-12, 
    4.318691e-12, 1.879275e-11, -5.998596e-13, -1.036324e-12,
  -2.512018e-13, -4.434092e-13, -4.794637e-13, -4.703876e-13, -4.539147e-13, 
    -3.792522e-13, -2.099709e-13, 1.229988e-13, 2.834677e-13, 4.697492e-13, 
    3.759493e-14, 4.642398e-13, 4.276579e-13, 8.110318e-13, 3.133327e-13, 
    -4.957562e-14, -1.711964e-14, -1.418032e-13, -5.320622e-13, 
    -3.055889e-13, -3.890638e-13, -9.91332e-13, -1.930428e-12, -7.580603e-13, 
    1.594697e-13, 1.060999e-12, -3.626266e-14, -3.388539e-13, -5.452028e-13, 
    -2.410849e-13, 1.64202e-13, 1.746797e-13, 7.771561e-13, -5.91055e-14, 
    -2.00992e-13, 4.463097e-14, -9.252543e-13, 5.108188e-13, -8.60978e-14, 
    -1.873487e-13, 5.221407e-13, -4.706652e-13, 1.4512e-13, -9.190131e-15, 
    -5.258294e-14, 3.948231e-14, -1.505088e-12, -7.853058e-13, 1.082162e-13, 
    1.576673e-13, -1.745753e-12, 1.343925e-13, 3.27452e-13, -6.756812e-12, 
    6.667819e-13, 4.19699e-13, -6.143419e-12, -2.140343e-13, -5.847601e-13, 
    2.371671e-12, -5.562079e-13, -5.388745e-13, 3.958778e-13, -1.196487e-13, 
    5.032086e-14, -7.272932e-13, -5.011269e-14, 4.066053e-13, 7.847056e-13, 
    2.144535e-13, -1.122713e-14, -2.964989e-13, 1.3059e-14, -1.899869e-13, 
    1.817726e-13, -1.447828e-12, -2.402523e-13, 1.240532e-12, -1.004835e-11, 
    -5.999368e-14, 7.915266e-13, -1.362372e-13, -9.756987e-13, 1.127182e-12, 
    6.702972e-14, -1.743466e-13, 3.053113e-16, -3.186201e-13, -6.160255e-13, 
    -8.609988e-13, -4.070771e-13, -2.132247e-12, 3.049436e-13, -3.218759e-13, 
    -2.262079e-15, -2.009636e-11, 1.233472e-12, 3.381045e-13, -3.992223e-12, 
    -1.730935e-12, 4.851952e-13, -1.909245e-13, 4.011808e-13, 7.153982e-13, 
    2.795125e-13, 2.03032e-13, 2.442768e-13, 5.805079e-14, -7.42878e-14, 
    1.12077e-13, 4.184986e-13, 1.4172e-13, 4.644896e-14, 1.722927e-13, 
    -2.156608e-14, 1.796317e-12, 5.476689e-12, 1.054812e-13, -2.320149e-13, 
    -2.070705e-13,
  -5.661166e-13, -3.402417e-13, -2.55726e-13, -3.524264e-13, -3.211181e-13, 
    -3.059358e-13, -2.790684e-13, 1.594141e-13, 4.034134e-13, -3.186201e-13, 
    5.219575e-13, 6.475237e-13, 5.192929e-13, 1.15602e-14, -3.835404e-13, 
    -1.674133e-13, -1.508377e-13, 6.505907e-14, -1.006244e-13, -6.120104e-15, 
    2.12011e-13, 3.51788e-13, -5.69364e-13, -4.278522e-14, 2.753214e-13, 
    2.740447e-13, 4.938411e-13, -3.118339e-14, -1.242478e-13, -1.802725e-14, 
    3.510109e-13, 5.816181e-14, -4.778816e-13, 8.034268e-13, -1.005598e-12, 
    2.970263e-13, -9.131945e-13, -4.52971e-14, -2.231951e-12, -2.957717e-13, 
    -8.426176e-13, -3.490402e-13, 8.715945e-14, 5.187257e-15, -3.279058e-12, 
    -2.004369e-13, -2.339795e-13, 4.286155e-14, -1.096293e-12, 2.065981e-11, 
    -2.62089e-13, -7.37424e-13, -1.40421e-13, -9.408336e-13, 4.597892e-13, 
    1.642367e-12, -4.279896e-12, -1.450828e-12, -2.422645e-13, 1.620502e-12, 
    9.505591e-13, -5.124096e-13, -6.123574e-13, -1.725758e-13, 1.132511e-13, 
    -4.234252e-13, 2.882833e-13, 1.507267e-13, 6.793177e-14, 3.965023e-13, 
    5.481032e-13, 4.028722e-14, -7.04839e-13, -3.755746e-13, 2.329664e-13, 
    -5.637574e-13, -2.115912e-13, -3.127082e-13, -4.088274e-12, 9.765799e-14, 
    6.755291e-13, 5.056178e-13, -1.249001e-16, -1.716266e-13, -7.100293e-13, 
    -1.180764e-12, 6.745993e-14, -3.554101e-14, -7.663817e-13, -4.131417e-13, 
    -1.714046e-13, 1.498354e-12, -3.783085e-14, 1.208569e-12, 6.916273e-13, 
    -3.433237e-12, -6.823708e-14, -4.476836e-13, 2.403119e-12, 3.019446e-13, 
    7.947393e-13, -1.739536e-12, 7.387788e-13, 3.379809e-12, -1.981887e-13, 
    1.393469e-13, 3.89952e-13, 8.69721e-14, -9.177381e-14, -4.601181e-13, 
    -6.139395e-13, -1.385433e-12, -5.463269e-13, -5.400264e-13, 3.60309e-13, 
    1.139641e-12, 3.540515e-12, -1.668277e-11, -1.724853e-12, -3.630568e-13,
  2.64927e-13, 1.499634e-13, -5.537237e-14, -1.143252e-13, 5.517808e-14, 
    4.650447e-13, 2.713108e-13, 3.420597e-13, 5.757061e-13, -7.426559e-13, 
    6.808443e-14, 7.019108e-13, 6.109002e-14, 4.536371e-13, -2.372158e-12, 
    -4.061584e-13, -6.549289e-13, 1.227074e-13, 3.748113e-13, 8.378853e-13, 
    2.03515e-12, -2.307876e-13, -2.254724e-12, -1.783296e-12, -7.91589e-13, 
    -3.031714e-12, -9.404144e-13, -5.705159e-13, -1.950023e-12, 1.105255e-12, 
    -3.01667e-12, -2.053996e-12, 6.73045e-13, -4.986289e-13, -1.432215e-12, 
    -8.666123e-13, -1.931261e-13, -3.21073e-13, -1.505879e-12, 7.165546e-13, 
    7.226553e-13, 1.642048e-12, -1.221176e-13, 7.77811e-14, -6.564888e-12, 
    1.196654e-12, 2.019218e-13, -9.058865e-13, -6.213363e-13, 3.101108e-11, 
    1.02756e-12, -1.146361e-12, 6.926376e-13, -3.376244e-12, 3.77641e-13, 
    1.30701e-13, 3.042289e-13, -7.703755e-13, 1.291744e-14, -7.814513e-13, 
    3.288869e-12, 2.417511e-14, 1.162404e-13, -7.28484e-13, -3.640532e-13, 
    -2.957301e-12, -1.590283e-12, 5.192791e-13, 1.32952e-12, -6.136203e-13, 
    -7.329692e-13, 2.642331e-12, -1.175199e-12, -4.671818e-13, 4.48111e-13, 
    -5.5983e-14, -3.027092e-14, -4.898582e-13, 2.984243e-12, 3.286427e-12, 
    1.539074e-12, 8.324897e-13, -8.830853e-13, -1.781908e-13, -1.15799e-12, 
    -5.2294e-12, -3.214207e-12, -2.084166e-13, 3.943742e-13, 1.240952e-13, 
    -1.377343e-12, 7.546131e-13, -1.165873e-13, 1.966533e-12, 2.329803e-12, 
    -1.208821e-11, -3.645195e-13, 1.988132e-13, 2.368103e-11, 1.679101e-13, 
    2.000927e-12, -8.411934e-13, 1.039949e-12, 4.233594e-12, -8.767986e-14, 
    -7.002732e-13, -1.206785e-12, -1.56189e-12, -8.106571e-13, -1.439654e-12, 
    -1.006223e-12, -1.532441e-12, -2.381428e-14, -8.731071e-13, 1.983996e-12, 
    1.243125e-12, 3.100541e-13, -4.693632e-12, -6.403645e-13, -2.02377e-12,
  6.311063e-13, 1.686429e-13, 5.932477e-13, 7.008283e-13, 2.547962e-14, 
    2.778888e-13, 2.678968e-13, 1.419087e-12, 6.542544e-13, 1.852074e-12, 
    5.909329e-12, 8.979595e-12, 7.94842e-12, 6.536161e-12, -9.389323e-12, 
    -1.736694e-12, 1.537714e-13, -2.009504e-13, -9.912904e-14, 1.640466e-12, 
    1.739997e-12, -6.455947e-13, -1.619704e-12, 3.151923e-13, -5.149381e-12, 
    -7.520429e-12, -3.387013e-12, -3.093636e-12, -4.832246e-13, 1.591838e-12, 
    -4.080181e-12, -3.980316e-12, 1.606271e-12, -2.424783e-12, -3.5838e-12, 
    -4.583389e-12, -2.243255e-12, -2.923356e-13, 5.984435e-12, 4.781731e-14, 
    -4.378497e-13, -6.374956e-12, 1.451436e-12, -1.4657e-12, -6.237066e-12, 
    7.989054e-12, 4.018452e-13, -2.790546e-13, 9.043877e-13, -1.90431e-13, 
    1.386717e-12, 1.97764e-12, -8.646806e-13, 4.872547e-12, -3.073569e-13, 
    -3.302081e-13, 4.302114e-14, 1.86251e-13, 6.908529e-13, 5.786427e-12, 
    -1.373845e-12, -1.277256e-12, -9.537371e-13, -5.835332e-13, 
    -1.409983e-13, -2.844613e-12, -6.012302e-12, 6.815715e-12, -7.784218e-12, 
    -1.145645e-11, -3.460232e-12, 3.926137e-12, -1.657563e-13, -7.231438e-13, 
    6.421141e-13, -1.681988e-14, -1.127015e-13, -2.810099e-12, -4.685155e-12, 
    7.561451e-12, 1.581263e-12, -3.955032e-12, 3.063105e-13, 2.134515e-12, 
    -3.469502e-12, -2.498057e-12, -9.181711e-12, -5.493384e-13, 
    -2.017683e-13, -1.39358e-12, -1.412537e-12, 7.90612e-13, -1.591505e-13, 
    1.470996e-12, 1.32111e-12, -3.823858e-12, 7.105982e-13, 9.535706e-13, 
    1.268563e-11, 2.541201e-12, 1.853628e-12, -1.458639e-12, 5.128918e-13, 
    4.466011e-13, 1.269596e-12, -1.373568e-12, -2.652212e-12, -2.48207e-12, 
    -1.001255e-12, -1.84619e-12, -1.255496e-12, -2.017275e-12, -2.381872e-12, 
    -2.545741e-12, -1.345407e-11, 4.254008e-12, 3.091263e-12, 1.674336e-12, 
    -9.971156e-13, -8.618661e-13,
  -4.375389e-13, -3.713252e-12, -2.443212e-12, -5.504097e-12, -4.513057e-12, 
    -4.541922e-12, -4.741818e-12, -5.181633e-12, 2.712713e-11, 2.471096e-11, 
    2.66403e-11, 1.197842e-11, 5.78515e-12, 6.492751e-12, -3.516742e-12, 
    9.821643e-13, -4.667994e-12, 1.411815e-12, 2.931787e-12, 1.213529e-12, 
    -1.565803e-12, -3.021194e-12, -2.711886e-12, -1.739331e-12, 
    -6.916911e-12, -5.001666e-12, -4.1675e-12, 2.529865e-12, 1.74199e-11, 
    -7.205347e-14, -2.008499e-11, 1.752914e-11, 2.533862e-12, 3.54583e-12, 
    -6.777856e-12, 1.338374e-12, -1.409195e-12, -3.942263e-13, -6.569023e-11, 
    -1.617317e-13, -2.694478e-12, -7.342515e-12, 3.394507e-14, 2.31884e-12, 
    2.098377e-12, -5.467515e-12, 1.619538e-13, 5.130063e-13, -2.739398e-12, 
    -1.119095e-11, 1.902228e-13, 1.02135e-12, 1.203926e-12, 1.529168e-11, 
    -2.665387e-12, -3.010647e-13, -5.137279e-12, 1.831535e-13, -7.805589e-13, 
    -1.166435e-12, 7.227552e-13, 4.427236e-12, -4.378276e-12, -5.884426e-12, 
    -6.118239e-12, 3.018386e-11, 2.013278e-11, -5.423884e-12, -8.305412e-12, 
    -1.347761e-11, -7.39192e-12, -1.394601e-11, 3.077927e-12, -2.770617e-12, 
    -1.991712e-12, -5.917489e-14, -7.244205e-15, 2.086248e-13, -7.524615e-12, 
    -2.881528e-12, -1.439643e-11, 6.637748e-12, -1.792622e-12, -1.027528e-11, 
    -2.821299e-12, 3.379075e-12, -3.815004e-12, 1.03334e-12, -8.820323e-13, 
    6.576406e-13, 2.330913e-13, -1.358239e-11, -1.229711e-13, 1.087225e-12, 
    1.312173e-12, -2.304657e-13, 2.407074e-13, 3.314182e-12, -3.291867e-12, 
    3.154144e-12, 4.849343e-12, -1.897173e-12, -2.178084e-13, -5.833747e-12, 
    -3.255063e-12, -8.223422e-13, -3.15703e-12, -3.933909e-12, -4.991452e-12, 
    -1.578626e-12, -3.535061e-12, -9.240775e-12, -3.305745e-12, 
    -5.261014e-12, -2.95125e-11, 1.008291e-11, 4.938536e-12, -5.316542e-12, 
    2.548656e-14, 9.426515e-12,
  -1.672207e-11, -2.920725e-11, -3.076983e-11, -2.21308e-11, -1.198697e-11, 
    -3.909206e-12, 4.72431e-11, 2.331219e-11, -5.568601e-12, -2.175488e-11, 
    -5.490552e-12, -1.466438e-12, -1.045386e-12, -1.593559e-12, 
    -1.280254e-12, -4.113376e-15, -7.96832e-12, 1.711048e-12, 4.131279e-13, 
    2.716716e-12, 4.21374e-12, 3.209044e-12, 7.600032e-13, 1.926348e-11, 
    5.361156e-12, 2.462336e-11, 2.536971e-12, 7.781498e-12, 1.710515e-11, 
    -1.247785e-11, -5.638934e-12, 1.191491e-12, 6.724343e-12, 8.410495e-13, 
    -2.607137e-12, 2.529532e-11, 3.225303e-12, -7.593648e-13, -8.162804e-11, 
    3.808065e-13, -1.350586e-13, -5.821288e-12, 4.455464e-12, 5.558129e-12, 
    -1.410816e-12, 1.055267e-12, -1.120021e-12, -7.830264e-13, 8.125045e-12, 
    -6.219286e-12, -1.176698e-12, -1.116218e-12, 8.685552e-13, 5.363487e-12, 
    -7.690889e-12, 5.769552e-13, -2.528866e-11, 2.81053e-13, -8.697932e-13, 
    -1.514201e-11, 2.476019e-12, 4.018008e-12, -2.559286e-12, -7.28344e-12, 
    -8.474887e-13, 7.637058e-12, 1.394124e-11, 4.854672e-12, 1.396494e-12, 
    4.061584e-12, 9.601209e-13, -1.89192e-11, 2.192135e-12, -2.912059e-12, 
    -2.724143e-12, 7.51621e-14, -1.494152e-13, -7.260942e-12, -1.062363e-11, 
    1.523892e-12, -2.790115e-11, 1.192388e-11, -3.238354e-12, -1.443901e-12, 
    -2.946754e-12, 2.190081e-12, -4.198641e-12, 1.968925e-12, 6.182051e-13, 
    3.688161e-13, 4.270362e-12, 5.769951e-12, 1.580402e-13, 2.92043e-12, 
    -7.919165e-12, 3.174128e-14, -2.524758e-12, -5.403289e-12, -1.108114e-11, 
    3.675449e-12, -8.546497e-13, -3.042809e-13, -7.715356e-14, -1.004711e-11, 
    -1.165179e-13, 1.758427e-12, 3.560374e-12, -5.210554e-12, -1.315292e-11, 
    9.005019e-13, -1.266282e-11, -2.5695e-12, -5.3203e-12, 2.025435e-12, 
    -1.40038e-12, 9.498046e-12, 2.148733e-12, -3.098362e-12, 7.023895e-13, 
    7.402634e-12,
  -5.561274e-12, 1.055059e-11, 1.663575e-11, 1.035461e-11, -8.001405e-12, 
    -4.311795e-11, 1.63575e-11, 3.099104e-12, -5.117998e-11, -1.356934e-11, 
    -5.654199e-12, -4.422157e-12, -2.706613e-12, 2.258221e-12, 2.938455e-12, 
    -3.512715e-12, -3.988906e-12, 3.874095e-12, 3.738055e-12, 4.013095e-12, 
    4.168998e-12, 3.026773e-12, 2.494172e-12, 2.70402e-11, 3.698375e-12, 
    -1.071088e-12, -1.257658e-11, 1.720291e-13, 1.311926e-11, -1.653466e-11, 
    -5.385281e-11, -1.21879e-10, -1.495903e-11, -9.775569e-12, -1.634692e-12, 
    -7.625539e-12, 3.812034e-13, -9.862146e-13, -7.999046e-11, -9.830192e-13, 
    -5.041667e-12, -5.836998e-12, 2.367662e-12, 5.676605e-13, 5.111828e-12, 
    3.395242e-11, -4.042183e-13, -1.626421e-12, 1.83206e-11, -1.322054e-12, 
    -1.186256e-12, -2.152145e-11, -6.093959e-13, -5.646039e-14, 
    -4.877087e-12, 5.509621e-13, -1.402931e-11, 5.633438e-13, -1.284312e-12, 
    -5.792922e-12, 6.680601e-12, -2.175898e-12, -2.255446e-12, -5.141259e-12, 
    -2.569123e-12, -4.188511e-12, -6.105993e-11, 8.426648e-12, 5.71912e-12, 
    -4.440556e-11, -1.029707e-11, -2.125883e-11, -3.344575e-12, 1.946851e-11, 
    -3.571393e-12, 8.34055e-14, -1.935327e-13, -5.559017e-11, -7.645205e-12, 
    -6.786238e-13, -2.565236e-11, 1.385379e-12, -1.538381e-12, -1.495143e-11, 
    -9.743345e-12, 7.046336e-12, -4.835882e-12, 5.060341e-12, 5.652458e-13, 
    -1.206396e-13, 7.576856e-12, -1.889022e-12, 1.227282e-12, -6.641596e-12, 
    -1.034123e-11, 1.845371e-12, 2.735034e-13, -1.329797e-11, -2.674583e-12, 
    3.34443e-12, -1.705691e-12, 7.285804e-13, 4.028652e-13, -4.81383e-12, 
    -6.329104e-12, 1.997874e-12, 1.138561e-12, 4.883455e-12, -1.111736e-11, 
    3.743283e-12, -2.14013e-11, 1.63613e-11, 1.907441e-11, 2.319647e-11, 
    6.721401e-12, -7.260747e-13, 1.81459e-13, -2.496178e-12, 5.279657e-12, 
    -1.513234e-12,
  1.360934e-11, 1.065942e-10, 4.095602e-11, -4.080047e-11, -8.690121e-11, 
    -4.525147e-11, -2.415923e-11, -2.413614e-11, -1.178696e-11, 1.256228e-11, 
    6.760537e-12, -3.662054e-11, -1.291334e-11, -8.641532e-12, -6.85918e-12, 
    -4.462925e-12, -4.652195e-12, 1.9032e-12, 4.984339e-12, 6.197043e-12, 
    6.045719e-12, 8.294032e-12, 6.964984e-12, 5.468459e-12, -1.452749e-11, 
    -2.49456e-11, -3.286982e-12, -1.495298e-11, 6.791734e-12, 1.279865e-12, 
    6.292117e-11, -9.506645e-11, -1.857242e-11, 7.769341e-13, -2.370149e-11, 
    -6.927015e-12, -1.641992e-12, -7.831513e-13, 1.143384e-10, -2.413658e-12, 
    -4.130718e-12, -1.919631e-11, 4.824099e-12, -1.219026e-12, 5.396794e-13, 
    7.478906e-12, 2.594314e-13, 1.776357e-14, 2.552924e-12, -2.821771e-13, 
    9.877807e-12, 3.704148e-12, -2.835615e-12, 9.873991e-13, 2.838854e-13, 
    4.571343e-13, -1.21127e-11, 9.269918e-13, -3.727274e-12, 9.580461e-12, 
    3.079759e-13, 1.646128e-12, -1.318501e-12, -9.313017e-12, -2.718203e-12, 
    -3.166356e-12, -1.31869e-10, 2.242095e-12, 8.593237e-12, -1.21692e-10, 
    -1.4172e-13, -4.239997e-11, -1.772044e-11, 1.649159e-11, -1.214862e-12, 
    -5.77316e-15, -2.549072e-13, 8.385972e-12, -1.033471e-12, -7.660539e-12, 
    -2.249045e-11, 1.366709e-12, 3.660933e-12, -2.895295e-11, -8.38396e-12, 
    2.128087e-11, -1.867367e-11, 1.619427e-12, -5.397245e-13, 3.670397e-13, 
    1.035666e-11, 3.956268e-12, 2.256223e-12, 1.088185e-12, -3.781975e-12, 
    6.307243e-12, 7.642109e-13, -2.84619e-11, 5.113687e-12, 9.01923e-13, 
    -2.525258e-12, 7.458881e-12, 3.62127e-13, -2.343764e-12, 1.35702e-11, 
    1.851824e-11, 5.700496e-12, 5.760503e-12, -1.325595e-11, -2.576828e-13, 
    -1.655515e-11, 2.635392e-11, 4.835105e-11, 1.353101e-11, 2.27568e-12, 
    -8.289591e-13, -8.900519e-14, -2.525931e-12, 5.762939e-12, -1.013012e-11,
  1.869119e-10, 6.981804e-11, -1.206601e-11, -7.11271e-11, -7.217593e-11, 
    -4.717049e-11, -5.557743e-11, -8.645784e-11, -4.13215e-11, -6.962997e-11, 
    4.460321e-12, -6.199707e-11, -7.027379e-12, -1.217282e-11, -5.731016e-11, 
    -4.568512e-12, -5.579737e-12, -2.132072e-12, 1.241449e-11, 4.992562e-12, 
    7.028378e-12, 5.241363e-12, 8.757217e-12, 4.02488e-11, -3.169931e-11, 
    3.618439e-12, -1.849765e-11, 1.006883e-11, 3.498091e-11, 5.606737e-11, 
    3.189704e-11, 1.051933e-10, -5.799516e-11, 1.232781e-11, -1.318301e-11, 
    4.225509e-12, 1.018907e-12, -2.311901e-13, 8.075707e-11, -4.271583e-13, 
    -6.409473e-12, -3.027401e-11, 3.101686e-12, -4.553562e-13, -7.088663e-12, 
    -8.01148e-12, 2.12963e-12, -9.777179e-13, 3.381517e-13, 1.698919e-13, 
    2.546151e-11, -9.617307e-12, -3.072054e-12, 1.0697e-12, 2.309575e-12, 
    3.898548e-13, -1.32927e-11, 1.256983e-12, 1.273981e-13, 1.32583e-11, 
    -6.461942e-12, 9.070522e-13, -4.670486e-12, -8.591062e-12, -3.546896e-12, 
    1.442135e-11, -2.556025e-10, 2.621836e-11, 4.296563e-12, -8.082202e-12, 
    2.204237e-11, 6.76843e-11, -4.800327e-11, -2.028455e-11, 8.944334e-12, 
    -7.893686e-14, 5.676015e-15, 3.064146e-11, 3.46062e-13, -6.545986e-12, 
    -1.774897e-11, 1.558034e-12, 2.225053e-12, -2.186795e-11, 4.773959e-15, 
    -1.152112e-11, -2.237688e-11, -7.545409e-12, -1.251122e-12, -4.20719e-13, 
    1.295908e-11, 3.177947e-12, 6.682987e-13, -3.557799e-12, -1.599965e-11, 
    7.539325e-12, 4.182965e-12, -6.797196e-11, 1.442935e-11, 3.110401e-13, 
    -2.237099e-11, 6.995231e-12, 4.462888e-13, -3.277933e-14, 5.588652e-11, 
    5.415135e-11, 3.992162e-11, 9.921841e-12, -1.60606e-11, -8.803513e-12, 
    -1.021083e-11, 2.784595e-11, 5.602474e-11, 9.248158e-12, -3.690381e-13, 
    -2.129963e-13, -2.054606e-13, -1.526324e-12, 2.169376e-12, 1.912581e-12,
  1.096492e-10, 7.641665e-12, -5.291545e-12, -3.832223e-11, -4.46978e-11, 
    -6.246714e-11, -8.094059e-11, -1.561817e-11, -9.006285e-11, -1.15278e-10, 
    -6.933654e-11, -3.847744e-11, -2.315992e-11, -7.505108e-14, 
    -1.115585e-10, -8.351475e-12, -5.744383e-12, 1.150602e-11, 8.021028e-12, 
    4.855227e-12, -1.675104e-12, -1.697309e-12, 1.733724e-11, 1.767009e-11, 
    9.064305e-12, -4.702683e-11, -3.044121e-11, 2.565237e-11, 5.523737e-11, 
    5.240275e-11, 1.981459e-11, 4.791323e-11, -6.893308e-11, -5.038303e-11, 
    4.543699e-12, -2.416534e-11, 1.780265e-12, 6.705747e-14, 2.70548e-11, 
    9.180434e-13, 3.537171e-12, -3.061196e-11, 7.072509e-12, 5.314811e-13, 
    3.285594e-12, 6.126655e-12, 5.187073e-12, -1.330491e-12, 6.439738e-13, 
    3.94268e-14, 3.96802e-12, -2.273892e-11, -8.005374e-13, 1.089884e-12, 
    5.344669e-13, 2.53908e-13, -2.265232e-11, 5.431877e-13, 1.990295e-11, 
    4.411138e-12, -9.063417e-12, -3.899348e-11, 3.348433e-12, -6.57856e-12, 
    -1.041212e-12, 9.267875e-11, -3.731726e-11, 3.520029e-11, 5.625722e-12, 
    5.110956e-11, 5.460765e-11, 2.143936e-10, -7.560841e-12, -2.594569e-11, 
    1.759906e-11, -2.833289e-13, 2.309541e-13, 2.5702e-11, 6.945833e-13, 
    -1.900347e-11, -1.661127e-11, -1.309791e-12, -2.702172e-12, 
    -8.121592e-11, 2.236056e-11, -6.595613e-12, -5.61919e-10, -1.279554e-11, 
    -8.737906e-13, -1.620926e-13, 4.681233e-11, 3.513945e-12, -6.271095e-13, 
    -2.390428e-11, -2.790457e-11, 5.895884e-12, 6.567991e-12, -7.565681e-11, 
    2.420109e-11, 1.186029e-12, -4.647127e-11, -1.35873e-11, 9.127837e-13, 
    1.738748e-13, 6.266143e-11, 2.518963e-11, 2.786571e-11, -4.544587e-12, 
    -1.732303e-11, -2.475353e-11, -1.246159e-11, 1.284617e-11, 5.849454e-11, 
    7.552847e-12, 6.253442e-12, 2.349454e-13, 3.885781e-16, -1.415326e-13, 
    6.737944e-13, 5.621725e-12,
  1.162515e-11, -4.638734e-12, -1.388645e-11, -4.899969e-11, -7.970535e-11, 
    -1.191178e-10, -1.380667e-10, -3.301648e-11, -1.712535e-10, 
    -2.972633e-10, -2.011677e-10, -9.866996e-12, -3.019784e-11, 2.773803e-11, 
    -5.359735e-11, -1.101523e-11, -4.057377e-12, 2.08813e-11, 1.246175e-11, 
    -4.298562e-12, -7.805978e-12, -2.402301e-12, 2.820344e-11, 8.34206e-11, 
    -9.139156e-11, -1.433718e-10, -3.247957e-11, 7.63849e-11, 1.223037e-10, 
    3.88114e-11, 8.439449e-11, 1.448315e-10, -5.224938e-10, -1.440708e-10, 
    -2.332687e-10, 4.611134e-11, -3.552269e-13, 2.359224e-13, 9.469692e-11, 
    -6.74838e-13, -2.33622e-12, -1.916667e-11, 5.899947e-12, 5.258849e-13, 
    -1.615954e-10, 2.565481e-11, 5.544232e-12, -3.499423e-13, 5.182077e-13, 
    -3.562706e-13, -1.666506e-11, 1.10203e-11, -5.519141e-13, 7.879475e-13, 
    -3.877898e-13, -1.654232e-13, -1.34172e-10, 5.20961e-13, 4.812906e-11, 
    -1.490108e-11, -3.160361e-12, -1.580707e-10, -1.510725e-11, 2.260281e-12, 
    2.19003e-11, -7.322492e-10, -8.563306e-11, 8.352008e-11, -8.679724e-13, 
    8.352496e-11, 1.875022e-10, 4.476102e-10, -4.067657e-11, -5.414846e-11, 
    9.742873e-12, -7.440715e-13, 7.127632e-14, 2.258616e-11, 1.135758e-14, 
    -1.097022e-10, -1.675327e-11, -9.641799e-12, -8.032686e-12, 
    -3.454903e-11, -4.46454e-11, -4.552401e-10, -2.866352e-11, -1.541722e-11, 
    -2.979422e-13, 3.876899e-13, 5.18654e-11, 2.96132e-12, -8.056888e-13, 
    -2.337024e-11, -4.536171e-11, 8.134826e-13, -3.288481e-13, 9.238454e-11, 
    2.647327e-11, 3.2363e-12, -2.622946e-11, 1.317494e-10, 7.75574e-13, 
    -7.64111e-14, 8.186629e-11, 3.259637e-11, 3.518408e-11, -1.06708e-11, 
    -3.20155e-11, -4.660472e-11, -2.271894e-11, -3.579137e-12, 3.889622e-11, 
    -5.67435e-12, 1.385447e-11, -5.706546e-14, 5.192513e-13, 1.22416e-13, 
    8.93452e-13, -4.344503e-11,
  2.913603e-11, -7.946976e-13, -4.384382e-11, -1.018214e-10, -1.486071e-10, 
    -1.851912e-10, -1.492457e-10, -4.225664e-11, -1.841538e-10, 
    -4.291942e-10, -4.192031e-10, -2.951903e-10, 3.565348e-11, 8.237877e-11, 
    1.509393e-11, -9.938939e-12, 2.055112e-12, 1.89877e-11, 2.285994e-11, 
    -3.443268e-11, -5.534906e-12, -4.634071e-13, 3.253686e-11, 6.424572e-11, 
    -5.715584e-11, -8.268564e-11, 1.705058e-11, 2.119951e-10, 2.214613e-10, 
    2.285394e-11, 1.667682e-10, 7.112377e-11, 4.491807e-11, -2.873255e-10, 
    -3.873166e-10, 2.452591e-10, -3.086287e-12, 1.960654e-13, 3.577985e-10, 
    -2.897105e-12, -3.708673e-11, 8.714141e-12, -7.78333e-12, -5.89459e-13, 
    -1.64311e-10, 1.469158e-11, 6.901368e-12, -4.980238e-12, 4.384493e-13, 
    -1.284306e-12, 1.530376e-11, -2.158163e-11, 2.97784e-12, 1.173328e-12, 
    9.280354e-13, -3.368417e-13, -4.513161e-10, 1.501954e-12, 5.138569e-11, 
    -2.470679e-11, 3.072431e-12, -2.804341e-10, -1.219262e-10, 2.272942e-11, 
    3.071503e-11, 3.906886e-10, 7.114598e-11, 1.620351e-10, 8.67062e-12, 
    1.288181e-10, 2.581511e-10, 5.715279e-10, 3.441543e-10, -7.76319e-11, 
    -1.319447e-11, -1.340927e-12, -1.164624e-13, 3.199085e-11, -1.493183e-12, 
    -2.154408e-10, -1.786726e-11, -1.473153e-11, -8.615553e-12, 
    -5.932743e-11, -5.249023e-11, -1.198905e-10, 1.553053e-10, -1.29512e-11, 
    -3.971823e-13, -3.318013e-12, 9.078271e-11, 3.582068e-12, -7.258638e-13, 
    -9.107337e-12, -8.071477e-11, -7.446621e-12, -1.4913e-11, -3.796585e-11, 
    2.648393e-11, 6.023493e-12, 2.100031e-11, 2.975197e-10, 7.588374e-13, 
    -1.972866e-13, 1.441782e-10, -5.876966e-11, 1.859157e-11, 1.627587e-13, 
    -3.618505e-11, -5.783529e-11, -3.070588e-11, -1.166156e-11, 
    -1.281419e-12, -3.368128e-11, 1.257949e-11, -2.247536e-13, 1.081357e-12, 
    -2.655653e-13, 2.117195e-13, -2.894864e-10,
  7.129675e-11, 1.046185e-11, -8.01208e-11, -1.689315e-10, -2.131033e-10, 
    -2.389537e-10, -1.511946e-10, -3.609646e-11, -5.145129e-11, 
    -1.124381e-10, -3.819061e-10, -7.553727e-10, 1.401776e-10, 1.467502e-10, 
    -7.827072e-11, -3.82574e-12, 3.288925e-12, 3.040368e-11, 2.044254e-11, 
    -6.262102e-11, -7.895018e-12, -4.620304e-12, 3.057998e-11, -6.39746e-11, 
    -2.007408e-10, -4.856746e-10, 2.206608e-10, 3.079901e-10, 2.833245e-10, 
    -5.382716e-11, 1.952891e-10, 1.789617e-10, 1.90342e-10, -2.031975e-11, 
    7.886225e-11, 3.774243e-10, -3.418687e-12, 2.4869e-14, 4.193774e-10, 
    -1.416236e-11, -4.367013e-11, 2.424283e-11, -1.888423e-11, -1.230488e-12, 
    -3.600853e-11, -1.434408e-12, 1.241451e-11, -3.28384e-11, 6.608047e-13, 
    -3.32534e-12, 5.936851e-11, -1.326237e-10, 2.890008e-11, 5.465495e-12, 
    3.56708e-12, 1.199041e-13, -5.204237e-10, 5.730438e-12, 3.785123e-11, 
    3.411527e-11, -7.503331e-12, -1.683897e-10, 2.265654e-11, 1.972236e-11, 
    1.862936e-11, 7.963319e-11, 8.175949e-11, 2.576783e-11, 3.321254e-11, 
    1.053531e-10, 2.28348e-10, 3.3081e-10, 1.073301e-10, -2.507061e-11, 
    -4.96005e-11, -2.499334e-12, 1.598721e-14, 3.483969e-11, 4.162226e-13, 
    -1.857661e-10, -2.034017e-11, -9.7371e-12, -1.885159e-12, 8.46816e-11, 
    -6.845813e-11, -3.240359e-10, 2.893872e-10, -7.233325e-12, -2.693054e-12, 
    -2.310774e-11, 5.441159e-11, 1.187978e-10, -2.144507e-12, 5.821565e-12, 
    -3.522871e-11, -1.926512e-11, -3.022098e-11, -2.395701e-10, 2.662581e-11, 
    7.435474e-12, -1.440448e-10, 1.218931e-10, 1.597722e-12, 3.167466e-13, 
    1.985496e-10, -3.173763e-10, -1.108758e-10, 2.30429e-11, -4.543654e-11, 
    -5.925749e-11, -3.553691e-11, -2.838174e-11, -4.632028e-11, 
    -6.316636e-11, 4.991563e-12, 3.552714e-15, 9.7089e-13, -4.964917e-13, 
    -1.96454e-12, -5.220437e-10,
  1.692566e-10, -1.886669e-11, -2.126637e-10, -2.399201e-10, -3.458744e-10, 
    -3.182645e-10, -2.212843e-10, -1.998224e-11, 3.508127e-11, 2.776925e-10, 
    -7.462297e-11, -2.524434e-10, 2.233076e-10, 1.898819e-10, -1.207905e-10, 
    7.600853e-12, 2.240341e-12, 5.069811e-11, 8.298473e-12, -7.018031e-11, 
    -1.37188e-11, -9.675816e-12, 1.722178e-11, -2.727951e-10, -5.286829e-10, 
    -8.59675e-10, -1.803802e-10, 3.201404e-10, -3.070184e-10, -2.055192e-10, 
    2.53646e-11, 4.51772e-10, 3.540901e-10, -1.044498e-10, 6.235332e-10, 
    4.890577e-10, -1.272227e-12, 1.316725e-13, 1.093525e-10, -5.443201e-11, 
    -2.032738e-10, 3.238299e-12, -1.440492e-11, -2.004313e-12, 4.230838e-10, 
    -4.196998e-11, 1.211653e-11, -1.492553e-10, 1.160316e-12, -6.691092e-12, 
    9.861534e-11, -2.804246e-10, 9.407462e-11, 1.017924e-11, 4.356959e-12, 
    3.321787e-13, -9.309673e-10, 1.200231e-11, 1.593623e-11, 2.686134e-10, 
    -2.214051e-11, 8.848033e-11, 1.617089e-10, 4.608936e-12, 2.10175e-11, 
    1.086526e-10, 1.817035e-11, -4.937171e-10, 7.938183e-11, 8.867218e-11, 
    2.491358e-10, -8.36188e-10, 2.476579e-10, 2.085372e-10, -6.541452e-11, 
    -4.474643e-12, 3.623768e-13, 1.892619e-11, 5.068657e-12, -1.047002e-10, 
    -3.019807e-11, 5.409007e-13, 1.090594e-11, -1.049649e-11, -7.251444e-11, 
    1.562352e-09, 4.032863e-11, 2.057376e-11, -1.398029e-11, -6.49063e-11, 
    7.038814e-11, 3.575632e-10, -1.538769e-12, 4.741292e-11, -1.971046e-11, 
    -3.000267e-11, -4.271961e-11, -4.188294e-10, 2.538059e-11, 7.894485e-12, 
    -5.283933e-10, -7.637102e-11, 2.979283e-12, -9.552359e-13, 1.657625e-10, 
    -3.608118e-10, -3.275833e-10, 1.421387e-10, -2.647127e-11, -5.249845e-11, 
    -2.900435e-11, -3.879208e-11, -7.396928e-11, -8.166801e-11, 
    -1.003109e-11, 9.256595e-13, -8.026912e-13, -1.846856e-13, -4.661493e-12, 
    -3.591953e-10,
  2.549481e-10, 2.52097e-10, -4.06791e-10, -5.708376e-10, -5.763425e-10, 
    -5.082992e-10, -4.44599e-10, 6.859757e-11, 4.930634e-11, -2.6332e-10, 
    -6.460805e-10, 3.645795e-11, 2.61382e-10, 2.351488e-10, -2.692957e-12, 
    2.472902e-11, 2.427036e-12, 5.474554e-11, 7.47602e-12, -6.205347e-11, 
    -1.811884e-11, -2.132694e-11, -6.034284e-12, -3.64464e-10, -8.328556e-10, 
    -1.068837e-09, -9.076953e-10, 9.208581e-10, -8.542145e-11, -3.312195e-10, 
    -8.812506e-12, 2.331326e-10, 1.882086e-10, 7.858247e-11, 1.111255e-09, 
    1.792539e-10, 1.396216e-12, 1.091127e-12, -6.250964e-10, -1.315604e-10, 
    -3.485546e-10, -4.340528e-11, -5.884182e-13, -2.155887e-12, 2.956853e-10, 
    -2.259686e-10, -8.07443e-12, -2.398015e-10, -3.722889e-12, -1.25352e-11, 
    2.072083e-10, -4.754401e-10, 1.125203e-10, 6.281909e-12, 8.473222e-13, 
    1.05782e-12, -5.38698e-10, 1.292175e-11, -3.559855e-11, 3.728409e-10, 
    -1.711165e-11, 2.118927e-10, 2.293241e-10, -3.521094e-12, 3.133422e-11, 
    -1.032543e-10, 4.066081e-12, -1.122338e-09, -2.440643e-10, 2.152571e-10, 
    4.712035e-10, -2.380933e-09, 1.506741e-10, 6.46553e-10, -3.629843e-11, 
    -5.545786e-12, 4.676259e-13, -1.599121e-11, 5.493606e-12, -1.001332e-11, 
    -5.764189e-11, -2.946962e-11, 2.64615e-11, 6.062706e-12, -3.460148e-10, 
    2.082826e-09, 3.108624e-13, 5.776357e-11, -4.458131e-11, -8.051071e-11, 
    4.545697e-11, 5.176354e-10, 7.232437e-12, 1.161814e-10, -1.828333e-10, 
    -2.715481e-11, -4.756373e-11, -6.059366e-10, 2.118483e-11, 6.620837e-12, 
    -4.852954e-10, -3.38384e-10, 2.971623e-12, -1.078104e-11, 1.097593e-10, 
    -7.362644e-11, -5.119745e-10, 1.942695e-10, -1.540243e-10, -6.375167e-11, 
    -1.658584e-11, -5.297807e-11, -1.019913e-10, -9.891643e-11, 
    -3.529799e-11, 2.99103e-12, -7.01661e-14, 4.45366e-13, -5.623835e-12, 
    -1.064393e-11,
  2.330864e-10, 4.753211e-10, 3.563976e-10, -3.058567e-10, -7.720757e-10, 
    -8.660734e-10, -7.821832e-10, 1.803038e-10, 1.443681e-10, 4.326779e-10, 
    -1.12307e-09, -2.331291e-11, 3.148735e-10, 3.415188e-10, 2.796021e-10, 
    3.949872e-11, 2.447287e-11, 2.924061e-11, 3.177369e-11, -4.600054e-11, 
    -2.793143e-11, -3.930367e-11, -2.509992e-11, -1.948841e-10, -1.42898e-09, 
    -1.66272e-09, -1.332232e-09, 1.553815e-09, -1.186006e-09, -4.234373e-10, 
    8.338219e-10, 3.273222e-10, 7.656205e-10, -4.007745e-10, 1.131156e-09, 
    -1.601492e-10, -2.001599e-12, 3.252509e-12, -1.437428e-09, -2.291028e-10, 
    -2.051593e-10, -1.490257e-10, 9.172219e-12, -2.312039e-13, -2.360075e-09, 
    -4.831833e-10, -1.464073e-11, -1.77101e-10, -1.368079e-11, -2.504796e-11, 
    1.076192e-10, 1.618616e-11, -1.462748e-10, -7.29301e-12, 2.184919e-12, 
    2.145839e-12, -1.040956e-09, 6.521006e-12, -3.948841e-11, -7.353411e-10, 
    3.318235e-11, 1.66164e-10, -8.304823e-11, -9.053025e-12, 3.055689e-11, 
    -9.689138e-10, -6.991101e-10, -9.124506e-10, -6.489849e-10, 4.397549e-10, 
    1.286768e-09, -2.614069e-09, -5.976837e-10, 1.472969e-09, -7.013093e-11, 
    -1.659117e-12, -1.807443e-13, -1.741274e-11, 6.702105e-12, -3.801404e-11, 
    -1.084892e-10, -7.954588e-11, 3.677236e-11, -6.028209e-10, -2.369163e-10, 
    8.362413e-10, 2.341061e-10, 9.653078e-11, -9.014295e-11, -1.521467e-10, 
    4.374066e-10, 2.779927e-10, 2.890665e-11, 1.62154e-10, -7.208172e-10, 
    -8.016698e-12, -4.805969e-11, -8.698429e-10, 1.751843e-11, -3.878853e-12, 
    -3.868266e-10, -4.723371e-10, -1.583178e-13, -3.162559e-11, 1.308678e-10, 
    2.369482e-10, -1.062244e-09, -1.115957e-09, -1.731042e-09, -5.084182e-10, 
    6.27054e-12, -6.451373e-11, -1.696208e-10, -2.05965e-10, -5.639222e-11, 
    6.708945e-12, 3.773426e-12, 1.583844e-12, -4.349188e-12, 2.088285e-10,
  2.14726e-10, 3.049365e-10, 5.185044e-10, 5.652296e-10, 3.000551e-10, 
    -3.751097e-10, -9.066738e-10, 1.386695e-10, 2.846363e-10, 6.262297e-10, 
    -8.870131e-10, -4.718004e-12, 3.282636e-10, 5.233147e-10, 7.843255e-10, 
    6.721734e-12, 5.478142e-11, 3.051781e-12, 4.851497e-11, -3.242917e-11, 
    -2.259526e-11, -4.519052e-11, -1.140421e-11, -2.005862e-11, 
    -2.611493e-09, -2.644114e-09, -1.698645e-09, 2.624532e-09, -8.02622e-10, 
    -2.986624e-10, 1.836554e-09, 1.306205e-09, 2.2291e-09, -7.836931e-10, 
    9.53257e-10, -6.514611e-10, 1.857074e-11, 6.199485e-12, -4.214229e-11, 
    -3.299618e-10, -2.37992e-10, -3.516405e-10, -9.610091e-13, 2.555511e-12, 
    -4.280899e-09, -6.168079e-10, 1.324167e-10, -1.691038e-10, -9.450218e-12, 
    -3.573453e-11, -4.728307e-11, 8.490062e-10, -5.780002e-10, -5.840804e-11, 
    5.043468e-11, 2.014389e-12, -4.11179e-09, 1.102975e-11, 1.87471e-10, 
    3.174998e-10, 1.062403e-10, 4.248335e-11, 3.737455e-10, -9.620749e-13, 
    1.89317e-11, -1.445933e-09, -3.513257e-09, 5.339373e-10, -7.709886e-10, 
    1.139121e-09, 2.265949e-09, -2.371017e-09, 3.103722e-10, 2.535586e-09, 
    2.58985e-10, 1.386979e-11, -1.499245e-12, 3.419487e-12, 2.99579e-11, 
    -1.202878e-10, -1.802043e-10, -1.72923e-10, 3.470291e-11, -1.678522e-09, 
    -1.202309e-10, -3.809774e-09, 4.070202e-10, 1.359695e-10, -1.138757e-10, 
    -3.51644e-10, 1.333873e-09, -3.02721e-10, 5.418066e-11, 1.515502e-10, 
    -2.194092e-09, 2.834355e-11, -6.183001e-11, -1.039552e-09, 1.712408e-11, 
    -2.248441e-11, 3.325624e-10, -8.510206e-10, -3.672174e-12, -6.593526e-11, 
    2.650822e-10, 3.469935e-10, -5.104823e-10, -2.03827e-09, -8.193695e-10, 
    -2.324661e-09, 5.046275e-11, -1.614353e-11, -3.530971e-10, -5.391669e-10, 
    -2.292211e-11, 1.173106e-11, 4.234835e-11, 3.006928e-12, -2.999823e-12, 
    2.002238e-10,
  1.530793e-10, 2.207088e-10, 6.100294e-10, 4.992842e-10, 7.77689e-10, 
    7.171366e-10, -3.492602e-10, -7.246115e-11, 1.47395e-10, 9.676313e-10, 
    -1.018449e-09, 2.195364e-09, 2.648335e-10, 7.337064e-10, 1.330761e-09, 
    -4.788347e-11, 7.035084e-11, 1.307399e-11, 4.228617e-11, -3.666401e-11, 
    -4.803269e-12, -1.814726e-11, 4.405365e-13, -5.621814e-11, -2.475119e-09, 
    -1.912753e-09, -1.80934e-09, 3.324573e-09, -4.483098e-10, -4.484946e-11, 
    2.314167e-09, 2.704425e-09, 2.126939e-09, -1.571266e-09, 9.04322e-10, 
    -1.062531e-09, 8.728165e-11, 9.359624e-12, -1.924533e-09, 1.583941e-11, 
    -5.198586e-10, -4.647802e-10, -3.917933e-11, -7.094325e-12, 
    -4.009905e-09, -5.579324e-10, 6.731469e-10, -3.023359e-11, 4.797585e-12, 
    -3.287504e-11, 9.370638e-11, 2.801244e-10, -6.59135e-10, -1.704308e-10, 
    1.009653e-10, -1.371347e-12, -3.001986e-09, 5.003358e-11, 3.419316e-10, 
    5.169909e-10, 1.490861e-10, -6.185985e-11, 8.263044e-10, 4.256435e-11, 
    3.552714e-11, -1.976261e-09, -4.030753e-09, 1.926892e-09, -3.644942e-09, 
    1.141927e-09, 1.141601e-09, -9.580958e-10, 3.53154e-10, 2.829893e-09, 
    1.972546e-09, 5.11875e-11, -3.755218e-12, -1.270379e-10, 7.57236e-11, 
    1.688392e-10, -2.695373e-10, -3.380027e-10, 5.2232e-11, -3.334577e-10, 
    -1.322746e-10, -3.600022e-09, 3.063718e-10, 1.672333e-10, -8.845724e-11, 
    -4.447998e-10, 1.77252e-09, -3.839261e-10, 7.912604e-11, 9.995915e-11, 
    -2.797776e-09, 7.020447e-11, -1.284917e-10, -8.334098e-10, 2.783906e-11, 
    -3.945786e-11, 4.630607e-10, -1.24401e-09, -5.432987e-12, -1.060751e-10, 
    2.892335e-10, 1.682565e-10, 5.884715e-10, 4.273915e-10, -5.670984e-10, 
    -2.149577e-09, -7.668177e-11, 7.261747e-11, -6.207159e-10, -1.025512e-09, 
    8.134293e-11, 1.202665e-11, 1.093401e-10, 2.881251e-12, -7.9039e-12, 
    8.689938e-11,
  3.074803e-10, -2.261331e-09, -4.3201e-11, 4.952483e-10, 3.979181e-10, 
    1.096069e-09, 4.553158e-10, -3.329035e-10, -3.895195e-10, 1.575629e-09, 
    -1.54067e-09, 1.708287e-09, 7.831744e-10, 1.045279e-09, 1.442061e-09, 
    -1.720991e-10, 1.602416e-11, 3.523581e-11, 6.78817e-11, -6.693313e-11, 
    1.483613e-11, 3.068124e-11, -7.7236e-11, -1.761748e-09, 1.013802e-09, 
    -1.096382e-09, -1.890186e-10, 4.832202e-09, 3.222524e-09, 1.105604e-10, 
    4.807632e-09, 2.876646e-09, 1.801425e-09, -1.690665e-09, 2.53678e-10, 
    -2.559645e-09, 3.106933e-10, 2.178702e-11, 3.806093e-10, 7.959472e-10, 
    -1.023346e-09, -2.930989e-10, -1.266898e-10, -6.048029e-11, 
    -4.214797e-09, -3.937259e-10, 1.607866e-09, -5.501022e-11, -4.222613e-11, 
    -7.831069e-12, 1.739195e-10, -6.615153e-11, 1.65852e-10, -2.010722e-10, 
    1.048747e-10, -8.149925e-12, 4.966125e-09, 1.304471e-10, 1.275504e-09, 
    3.926486e-09, 9.065104e-11, -1.842864e-10, 1.976304e-10, 1.980766e-10, 
    9.155485e-11, -5.26947e-09, -6.581985e-09, -1.887145e-09, 1.477574e-09, 
    3.082434e-09, -1.538936e-09, 2.343512e-10, 4.15767e-10, 1.740787e-09, 
    2.794901e-09, 8.176926e-11, -7.029044e-12, -4.06164e-10, 3.405383e-11, 
    1.382759e-09, -3.575735e-10, -6.028852e-10, 1.637801e-10, -4.161791e-10, 
    -3.82741e-10, 5.492211e-10, 3.531255e-10, 1.644338e-10, -1.090199e-10, 
    -1.141807e-09, 1.324963e-09, 6.559446e-10, 9.611867e-11, 1.527098e-10, 
    -2.817401e-09, 9.614922e-11, -2.768132e-10, -7.494378e-10, 6.474465e-11, 
    -7.585754e-11, 4.247624e-10, -1.576651e-09, -9.778844e-12, -1.44043e-10, 
    2.208367e-10, -1.506208e-10, 3.928022e-10, -6.456986e-10, -2.379295e-09, 
    -9.909229e-10, -5.66061e-10, 8.550671e-11, -9.464287e-10, -1.231186e-09, 
    2.061569e-10, 1.490292e-11, 1.0359e-10, -6.277201e-12, -2.826628e-11, 
    3.871037e-11,
  9.328005e-10, -6.194796e-10, -5.233403e-09, -2.242444e-09, -1.129422e-09, 
    3.407195e-10, 1.590507e-09, -8.786571e-11, -1.245397e-09, 2.100236e-09, 
    3.957581e-10, -2.267072e-09, 1.646995e-09, -6.52193e-10, 9.042793e-10, 
    -5.836497e-10, -3.148017e-10, -9.80549e-12, 1.694307e-10, -3.497291e-11, 
    4.874323e-12, 1.271871e-11, -1.863754e-10, -2.760601e-09, 5.946987e-09, 
    3.786909e-10, -3.414158e-10, 7.299576e-09, 1.090685e-08, -3.288818e-10, 
    -1.109726e-09, 1.267239e-09, 1.304684e-09, -6.248655e-10, -4.174723e-10, 
    -4.786941e-09, 6.723397e-10, 4.753709e-11, 6.083795e-09, 1.294173e-09, 
    -1.76754e-09, -5.388756e-11, -5.650378e-10, -1.759175e-10, -7.721965e-09, 
    -3.287681e-10, 2.736442e-09, -8.348877e-12, -5.196398e-10, 3.519229e-11, 
    1.593463e-10, 4.75211e-11, 4.171241e-10, -1.991822e-10, 2.066184e-10, 
    -1.394085e-11, 2.003432e-08, 2.483077e-10, 1.100493e-09, -1.04234e-09, 
    -8.839152e-12, -4.87546e-10, -1.1255e-11, 1.441899e-09, 7.994742e-11, 
    -1.018981e-08, -3.175714e-09, -2.173948e-09, 7.500205e-10, 2.821409e-09, 
    -2.368353e-09, 1.148791e-09, 5.163798e-10, 1.721403e-09, 3.371086e-09, 
    6.241407e-11, -6.082246e-12, -6.773249e-10, -1.896076e-10, 1.677037e-09, 
    -4.021246e-10, -1.036287e-09, 4.373888e-10, 2.719645e-09, -2.506226e-10, 
    8.135004e-10, 1.035147e-09, 1.353442e-10, -1.81686e-10, -1.820325e-09, 
    7.105712e-10, 1.311855e-09, 1.006768e-10, 2.182304e-10, -2.57559e-09, 
    1.229239e-10, -4.560036e-10, -1.043887e-09, 1.324736e-10, -1.234753e-10, 
    -1.499671e-10, -1.751684e-09, -2.026646e-11, -1.5888e-10, 1.378169e-10, 
    -5.52177e-10, -2.898304e-10, -1.282899e-09, -2.591349e-10, -3.141821e-09, 
    4.29722e-10, -1.849401e-10, -9.666934e-10, -1.118408e-09, 3.584262e-10, 
    1.771525e-11, -2.134275e-10, -2.825207e-11, -6.467449e-11, -1.976446e-10,
  2.242022e-09, -2.328616e-09, 2.092978e-09, -5.312923e-09, -7.025303e-09, 
    -5.084893e-10, 1.974772e-09, 1.03859e-09, -2.933653e-10, 2.966377e-09, 
    6.009973e-09, -2.960316e-09, 2.82532e-09, 1.783523e-09, -9.822188e-11, 
    -8.79421e-10, -6.828422e-10, -4.646061e-10, 3.988134e-10, 5.11946e-12, 
    -3.424461e-11, -5.672618e-11, -1.338343e-10, -2.19887e-09, 9.672394e-09, 
    5.513531e-09, 1.013749e-09, 1.083081e-08, 1.184114e-08, 2.643574e-11, 
    -4.139022e-09, 4.985523e-11, 3.365674e-09, -1.720249e-09, -7.774155e-10, 
    -6.372343e-09, 9.914466e-10, 7.147349e-11, 9.025886e-09, 9.984582e-10, 
    -2.50973e-09, -9.560708e-11, -1.469903e-09, -4.075393e-10, -6.790682e-09, 
    8.708767e-11, 4.251678e-09, 1.649987e-10, -8.867992e-10, 7.458922e-12, 
    1.04329e-10, -8.978382e-10, 7.39832e-10, 1.445734e-10, 2.122292e-10, 
    -1.31557e-11, 3.121139e-08, 4.030149e-10, 1.271852e-09, -7.760903e-10, 
    -6.411582e-11, -7.519212e-10, -5.962519e-11, 4.271451e-09, 4.152199e-11, 
    -1.606747e-08, 3.08933e-09, -4.673151e-09, -5.86536e-09, 2.370431e-09, 
    -3.222702e-10, 4.238533e-09, 8.181793e-10, 1.735916e-09, 2.803896e-09, 
    4.780887e-11, 1.196199e-11, -7.189307e-10, -2.627445e-11, 1.596479e-09, 
    -8.127294e-10, -1.685306e-09, 8.570034e-10, 4.88328e-09, 1.019121e-09, 
    5.341896e-10, 1.266333e-09, 1.348646e-10, -2.012035e-10, -3.044445e-09, 
    -1.053273e-10, 1.292663e-09, 9.596945e-11, 8.666419e-11, -2.003528e-09, 
    1.811749e-10, -5.290211e-10, -5.115588e-10, 2.033893e-10, -1.805141e-10, 
    -6.870913e-10, -1.688107e-09, -4.557599e-11, -1.123865e-10, -1.37387e-10, 
    -1.48469e-09, -1.946827e-09, -3.074344e-09, -3.874501e-09, 7.580425e-11, 
    3.2278e-09, 8.123813e-10, -1.157101e-09, -8.003802e-10, 6.860752e-10, 
    -7.519674e-12, -4.726388e-10, -4.339906e-11, -9.653789e-11, -5.09683e-10,
  4.286012e-09, 1.081151e-09, -5.062855e-09, -6.247557e-09, -9.414503e-09, 
    -5.135075e-09, 1.300652e-09, 2.972104e-09, 1.806615e-09, 3.566658e-09, 
    7.495903e-09, 2.994955e-09, 3.090936e-09, 4.288172e-09, -9.501484e-10, 
    -9.665704e-10, -6.42941e-10, -1.026674e-09, 1.22942e-09, -1.155581e-09, 
    -7.407763e-11, -3.034977e-10, 2.392042e-11, -3.308394e-10, 1.11706e-08, 
    7.912224e-09, 2.344553e-09, 1.300949e-08, 1.240081e-08, 1.885457e-09, 
    5.861871e-10, 5.785701e-10, 1.763755e-09, -4.296293e-09, -4.687983e-10, 
    -6.506252e-09, 1.193843e-09, -9.841017e-13, 7.583356e-09, 7.86526e-10, 
    -3.434729e-09, -6.94552e-10, -1.494126e-09, -6.915188e-10, -2.314192e-09, 
    3.81835e-10, 8.904397e-09, 2.753247e-10, 9.726542e-11, -1.138396e-10, 
    -1.279084e-10, -2.62413e-09, 1.06993e-09, -8.348522e-11, 1.842743e-10, 
    -1.071143e-11, 2.605536e-08, 6.104877e-10, 6.089235e-09, -2.68443e-10, 
    4.176925e-11, -6.776695e-10, -5.255565e-10, 4.704044e-09, 1.476231e-10, 
    -2.207225e-08, 2.658954e-09, -5.273858e-09, -1.953852e-08, 2.313175e-09, 
    5.073737e-10, 7.58563e-09, 1.190376e-09, 1.415277e-09, -9.344653e-10, 
    8.812506e-11, 2.632561e-11, -6.726388e-10, 9.751062e-11, 8.388561e-10, 
    -2.646711e-09, -2.275128e-09, 1.48454e-09, 2.433655e-09, -9.887451e-10, 
    -6.055636e-10, 4.767635e-10, 1.912106e-10, -2.02574e-10, -2.886363e-09, 
    -2.478071e-09, 1.944142e-09, 7.105072e-11, -3.078292e-10, -4.873009e-10, 
    2.676849e-10, -4.533199e-10, 1.848083e-09, 2.513794e-10, -2.463246e-10, 
    -5.016823e-10, -1.367635e-09, -1.01025e-10, -2.530776e-11, -8.757119e-10, 
    -1.918504e-09, -2.686516e-09, -6.195688e-09, -6.569518e-09, 9.93527e-10, 
    6.634327e-09, 6.60453e-10, -1.439854e-09, -5.151541e-10, 1.344933e-09, 
    -4.017622e-11, -2.84551e-10, -2.593037e-11, -1.065086e-10, -6.507825e-10,
  5.958356e-09, -2.674767e-09, -7.696485e-09, -5.793112e-09, -1.770275e-09, 
    -1.006708e-08, 1.250129e-09, 3.711449e-09, 2.173095e-09, 4.204225e-09, 
    9.427652e-09, 8.089046e-09, 4.591612e-09, 2.019249e-09, -1.363617e-09, 
    9.473222e-11, -3.698943e-10, -1.420617e-09, 3.411287e-09, -7.17165e-10, 
    -1.186606e-10, -6.828316e-10, 1.707576e-10, 1.170207e-09, 1.158088e-08, 
    6.138777e-09, 2.232724e-09, 1.339481e-08, 9.487024e-09, -4.477272e-09, 
    2.545363e-09, 3.4305e-11, 2.761738e-09, -7.048357e-09, -2.195577e-10, 
    -7.394249e-09, 1.119025e-09, -1.926423e-10, 8.396626e-10, 1.336304e-10, 
    -3.020801e-09, -7.59627e-10, 1.345768e-11, -8.699161e-10, 2.739142e-09, 
    1.364157e-09, 2.19882e-08, 3.6394e-11, -6.154834e-10, -1.677822e-10, 
    -4.188756e-10, -3.188575e-09, 1.419048e-09, -1.310013e-10, 4.819185e-10, 
    -2.184208e-11, 3.137521e-08, 8.905715e-10, 1.931924e-08, 6.119194e-11, 
    3.269065e-10, -1.115268e-09, -1.044043e-09, 2.071827e-10, 4.062997e-10, 
    -2.481875e-08, -1.076046e-10, -2.263022e-09, -2.52177e-08, 4.476988e-10, 
    -4.429239e-10, 9.311634e-09, 4.3309e-10, -4.405365e-11, 6.861797e-10, 
    8.901679e-11, 2.576428e-11, -1.066191e-09, 2.721343e-10, 8.333245e-10, 
    -4.850108e-09, -2.697274e-09, 2.290562e-09, -2.79357e-10, 1.60523e-09, 
    -4.590959e-10, 6.755556e-10, 2.258673e-10, -4.270455e-10, -1.239556e-09, 
    -9.334343e-09, 3.674444e-09, -3.304024e-11, 7.235343e-10, -5.582592e-10, 
    3.490726e-10, -3.734158e-10, 4.793264e-09, 3.378773e-10, -3.641787e-10, 
    -6.122036e-11, -2.021277e-09, -2.233858e-10, 1.200107e-11, -1.130815e-09, 
    -1.096879e-09, -2.641855e-09, -7.880885e-09, -5.995958e-09, 1.209912e-09, 
    1.281367e-08, 2.491447e-10, -2.258815e-09, -4.912692e-10, 1.694019e-09, 
    -2.237641e-11, -1.014335e-10, 2.356959e-11, -9.852918e-11, -6.816663e-10,
  5.726292e-09, -7.55108e-10, -8.873826e-10, -2.889522e-09, 8.241727e-10, 
    -6.468667e-09, 8.541292e-10, 4.383594e-09, 1.819046e-09, 4.460219e-09, 
    6.737821e-09, 1.721327e-08, 5.263871e-09, -5.582592e-10, 2.43233e-10, 
    -8.265659e-10, -2.788056e-10, -1.876401e-09, 6.488548e-09, 1.137039e-09, 
    -2.852971e-10, -8.954544e-10, 1.201101e-10, 5.867378e-10, 6.070763e-09, 
    7.841095e-09, 1.989292e-09, 1.270331e-08, 3.50833e-08, -1.025631e-08, 
    7.047163e-09, 6.235723e-11, 6.434902e-09, -9.498365e-09, 3.919922e-10, 
    -8.618258e-09, 2.494119e-10, -2.70802e-10, -3.535547e-09, -4.839533e-10, 
    -1.362685e-09, -1.193143e-10, 1.798654e-09, -1.241153e-09, -1.175238e-09, 
    2.992806e-09, 3.824357e-08, 3.051355e-10, -1.767762e-09, -1.726441e-10, 
    -6.900152e-10, -1.105263e-09, 2.763613e-09, -4.241997e-10, 4.046555e-10, 
    -4.541789e-11, 4.328086e-08, 1.131298e-09, 2.822254e-08, -4.912692e-11, 
    4.485514e-10, -2.50418e-09, -1.416709e-09, -7.359995e-09, -1.38823e-10, 
    -1.755586e-08, -6.209177e-09, 2.754348e-09, 4.0896e-09, 4.856645e-09, 
    -9.657697e-10, 7.444328e-09, 1.972467e-11, -1.18257e-09, 9.920598e-10, 
    8.526513e-12, 1.337952e-11, -2.195321e-09, 5.32404e-10, 1.520391e-09, 
    -5.262848e-09, -3.722523e-09, 3.200682e-09, -1.300918e-09, 7.884751e-10, 
    -4.461072e-10, 1.967408e-09, 2.331149e-10, -1.212402e-09, 3.545608e-10, 
    -1.141922e-08, 5.405855e-09, -1.774509e-10, 6.64636e-10, 2.783054e-10, 
    4.963908e-10, -4.525305e-10, 6.845369e-09, 4.992557e-10, -4.766548e-10, 
    3.438686e-09, -5.236739e-09, -4.396341e-10, -6.846435e-11, -4.607159e-10, 
    -3.688001e-10, -1.920682e-09, -2.732975e-09, -2.764182e-09, 4.770527e-09, 
    1.945421e-08, -1.062574e-09, -4.050491e-09, -5.68491e-10, 4.589538e-10, 
    -4.956746e-12, -3.67848e-11, 8.776446e-11, -9.636025e-11, -4.264393e-10,
  3.573405e-09, 3.773266e-10, 9.820269e-10, 4.99881e-10, 2.462457e-10, 
    7.154881e-10, -2.613604e-09, 4.365859e-09, 3.480068e-09, 2.214392e-09, 
    4.660876e-09, 1.336315e-08, 4.528886e-09, 1.011131e-09, 2.409479e-09, 
    -2.137779e-09, -4.042135e-11, -2.665644e-09, 8.663292e-09, 2.031982e-09, 
    -2.153342e-09, -9.730456e-10, -1.098783e-10, -5.186394e-10, 1.201499e-09, 
    9.367739e-09, 2.746333e-09, 2.380716e-09, 1.858029e-08, -1.652131e-08, 
    6.215146e-09, -2.831939e-10, 1.000001e-08, -8.970801e-09, -2.974048e-10, 
    -9.248083e-09, 1.020339e-10, -4.848033e-11, -2.735703e-09, -1.102372e-10, 
    1.825936e-09, 6.136816e-10, 3.597293e-09, -1.377115e-09, -1.148635e-09, 
    6.947573e-09, 3.807165e-08, 1.723123e-09, -3.425168e-09, -2.51724e-10, 
    -6.990817e-10, -6.796199e-10, 3.999378e-09, -1.855483e-10, -3.344112e-10, 
    -2.751221e-11, 5.032763e-08, 1.021982e-09, 2.356355e-08, -1.666464e-09, 
    -2.904699e-11, -2.919649e-09, -1.765329e-09, -9.446353e-09, 
    -4.072945e-09, -2.362356e-09, -8.30272e-09, 1.238851e-08, 2.166303e-09, 
    9.174414e-09, -1.812168e-10, 2.505658e-09, -2.634692e-10, -2.227694e-10, 
    -2.788971e-09, -5.815082e-11, 4.263256e-12, -3.944322e-09, 9.250911e-10, 
    4.113872e-09, -5.442587e-09, -6.337314e-09, 3.872714e-09, 3.529237e-09, 
    -3.413049e-09, 1.997194e-09, 2.564832e-09, 1.894023e-10, -1.695672e-09, 
    6.62169e-10, -1.906415e-09, 7.70866e-09, -7.076579e-10, -9.865857e-09, 
    4.182141e-09, 1.280705e-09, -6.811434e-10, 6.086282e-09, 5.152287e-10, 
    -5.621814e-10, 3.358707e-09, -5.77516e-09, -5.736425e-10, -3.197513e-10, 
    3.618084e-10, 1.875264e-10, -5.287006e-10, 2.803517e-10, -2.417266e-09, 
    9.091366e-09, 1.580293e-08, -1.43848e-09, -7.181313e-09, -3.503828e-10, 
    -1.094691e-09, -2.411298e-11, 9.469403e-11, 1.39277e-10, -1.029896e-10, 
    2.214051e-10,
  1.250328e-09, 1.756973e-09, -3.933565e-11, 3.750529e-10, -9.840733e-10, 
    2.50003e-09, -9.338862e-09, 3.178059e-09, 5.62062e-09, -1.017384e-09, 
    3.58807e-09, 8.02271e-09, -4.63217e-10, 1.120702e-08, 7.022663e-09, 
    -1.216153e-09, -4.420144e-11, -1.379135e-09, 9.720175e-09, 6.702749e-09, 
    -7.075244e-09, -1.199567e-09, -1.259252e-09, -1.713943e-09, 
    -4.263256e-11, -2.442562e-10, 4.208232e-09, 8.231552e-09, -2.875822e-09, 
    -1.280932e-08, 2.787431e-09, -1.950355e-09, 1.363327e-08, -1.049602e-08, 
    -4.975789e-09, -1.05141e-08, -5.535014e-10, 2.498268e-10, 1.444732e-09, 
    1.015094e-09, 5.951676e-09, 1.652438e-10, 4.169664e-09, -1.463544e-09, 
    -6.157336e-09, 1.376054e-08, 3.51437e-08, 3.254002e-09, -5.229549e-09, 
    -3.26537e-10, -4.978133e-10, 1.161141e-09, 4.450436e-09, -2.743832e-10, 
    1.111866e-09, 5.275069e-11, 4.909532e-08, 6.203607e-10, -1.281784e-08, 
    -6.24199e-09, -3.942375e-09, -2.454669e-09, -8.66919e-10, -9.098085e-09, 
    -8.68589e-09, 1.013927e-08, -7.341498e-09, 3.120482e-08, 1.449848e-09, 
    7.073083e-09, 3.523155e-10, 1.408068e-09, -2.335696e-10, 8.390089e-11, 
    -2.435593e-09, -4.888534e-11, -1.128768e-10, -6.299771e-09, 1.505225e-09, 
    5.249944e-09, -6.1994e-09, -1.057915e-08, 3.731827e-09, 4.195954e-09, 
    -3.205741e-09, 1.121691e-09, 1.335309e-09, 1.442118e-10, -4.422504e-09, 
    -3.995524e-10, 1.325708e-08, 1.188773e-08, -2.097394e-09, -1.483076e-08, 
    6.523067e-09, 4.236762e-09, -9.646215e-10, -6.787673e-10, 4.081926e-10, 
    -7.934546e-10, 1.657213e-09, -1.578542e-10, -3.939711e-10, -6.586696e-10, 
    2.630316e-09, 1.462013e-09, -7.889298e-10, -1.757996e-09, -4.846754e-09, 
    7.762253e-09, 8.279983e-09, -5.453558e-10, -1.031771e-08, 2.323191e-10, 
    2.863771e-10, -7.599965e-11, 2.61025e-10, 1.621476e-10, -1.146034e-10, 
    -8.520828e-11,
  -5.894663e-11, 1.595879e-09, -1.425178e-09, -1.094918e-09, -1.48674e-09, 
    -7.778453e-10, -1.411507e-08, 2.753325e-09, 4.880633e-09, -6.559731e-10, 
    2.307843e-10, 5.17889e-09, -1.125312e-08, 1.005662e-08, 7.557105e-09, 
    -2.62528e-09, -7.021811e-10, -3.108198e-10, 9.829066e-09, 1.230438e-08, 
    -9.656276e-09, -1.208321e-09, -3.033961e-09, -3.100524e-09, 
    -7.101448e-10, -1.323201e-09, 1.651921e-08, -1.197839e-08, -8.738482e-09, 
    -1.507829e-09, -2.779359e-09, -4.8571e-09, 1.841312e-08, -1.326379e-08, 
    -4.487504e-09, -1.330312e-08, -5.108063e-10, 5.440484e-10, -2.716149e-09, 
    2.985972e-09, 1.072551e-08, -1.034874e-08, 9.724502e-09, -7.684227e-10, 
    -2.881222e-09, 1.874946e-08, 4.032847e-08, 3.735138e-09, -5.507093e-09, 
    -4.00135e-10, 1.329425e-11, 2.441425e-09, 5.356083e-09, -3.971422e-10, 
    4.30731e-09, 1.844285e-10, 3.187762e-08, 8.113034e-10, -1.056877e-08, 
    -1.287662e-08, -1.081821e-08, -1.402043e-09, 3.524292e-12, -1.317237e-08, 
    -5.026731e-09, 3.159244e-09, -9.677024e-10, 4.292394e-08, 1.56337e-08, 
    -4.140304e-09, -4.592948e-10, 1.532391e-08, 6.061782e-10, -3.47768e-10, 
    7.269647e-10, 4.092726e-11, -2.073008e-10, -1.03791e-08, 2.406892e-09, 
    -7.827566e-09, -1.075475e-08, -1.583967e-08, 2.632078e-09, 1.124306e-09, 
    1.235207e-09, 2.455522e-09, -1.175977e-09, -8.969891e-11, -7.605194e-09, 
    -3.299675e-09, 1.308433e-08, 2.0877e-08, -4.371771e-09, -2.936991e-08, 
    6.497828e-09, 9.656446e-09, -1.224748e-09, -7.261178e-09, -4.453113e-10, 
    -1.260878e-09, 2.177671e-10, 2.119574e-09, 6.436451e-11, -1.091024e-09, 
    1.022386e-08, 5.017341e-09, 2.42278e-09, -8.825225e-09, -4.573337e-09, 
    5.871641e-09, 3.000309e-09, -6.288019e-10, -7.184724e-09, 1.351566e-09, 
    2.106333e-09, -1.855028e-10, 4.505054e-10, 2.080345e-10, -8.984102e-11, 
    -1.420233e-09,
  9.487167e-11, 2.008278e-10, -2.140951e-09, -1.422165e-09, -1.548472e-09, 
    -2.456602e-09, -1.087858e-08, 3.203525e-09, 4.757794e-09, 2.084391e-09, 
    -3.462333e-09, 1.512262e-09, -1.298827e-08, -1.498847e-09, 7.535846e-09, 
    -2.950792e-09, -1.110533e-09, 6.72884e-10, 8.523884e-09, 1.371467e-08, 
    -5.58174e-09, -4.16486e-09, -4.333856e-09, -1.804324e-09, -5.038601e-10, 
    5.950938e-10, 2.779882e-08, -3.061444e-08, -2.623722e-09, 1.234997e-08, 
    -6.692176e-09, -7.797041e-09, 2.090798e-08, -1.601103e-08, -5.08976e-10, 
    -1.648232e-08, -1.146122e-09, 9.215455e-10, -1.272383e-08, 3.793183e-09, 
    1.69092e-08, -1.55228e-08, 1.294434e-08, 3.010481e-10, -6.770676e-09, 
    3.164928e-09, 4.914369e-08, 4.437766e-09, -6.509435e-09, -6.483099e-10, 
    1.233232e-09, -1.029264e-09, 8.306097e-09, -5.392394e-10, 2.377763e-09, 
    3.334435e-10, 6.945385e-08, 3.631516e-09, 8.908896e-10, -1.877328e-08, 
    -9.355119e-09, 3.411742e-09, 1.228386e-10, -1.877637e-08, 8.106213e-10, 
    -3.53748e-09, 4.678157e-09, 3.816052e-08, 9.39832e-09, -3.484217e-09, 
    -1.767319e-09, 2.570715e-08, -2.820116e-09, -1.087699e-09, 9.002838e-09, 
    1.513172e-10, -9.829648e-11, -1.745309e-08, 3.58268e-09, 2.27999e-09, 
    -1.629559e-08, -1.991162e-08, 8.918164e-10, 3.883542e-10, 6.84912e-09, 
    4.362164e-09, -2.126399e-09, -1.233161e-09, -9.886682e-09, -9.25769e-09, 
    6.136361e-09, 3.002546e-08, -5.560324e-09, -2.696239e-08, 7.370261e-09, 
    1.661899e-08, -1.495948e-09, -2.846502e-08, -2.297782e-09, -2.167963e-09, 
    -1.03114e-09, 7.223896e-09, 3.046132e-10, -1.376506e-09, 1.276288e-08, 
    7.653057e-09, 4.843059e-09, -2.059983e-08, 2.08081e-09, 5.877894e-09, 
    2.752188e-09, -2.826198e-09, 1.257661e-09, 2.167042e-09, -8.808456e-10, 
    -3.873879e-10, 6.89802e-10, 2.730935e-10, -4.147083e-11, -3.169305e-09,
  1.231399e-09, -8.491838e-10, -2.682839e-09, -9.122232e-10, -4.922072e-10, 
    -1.841784e-09, -7.959216e-10, 1.578428e-09, 8.256109e-09, 3.819764e-09, 
    -2.301022e-09, 7.497647e-11, -9.748874e-09, -9.614723e-09, 1.710725e-08, 
    -3.841187e-09, -3.666849e-09, 6.687628e-11, 6.458677e-09, 9.108305e-09, 
    8.503775e-10, -9.0605e-09, -3.72529e-09, 4.334652e-09, 4.078515e-10, 
    1.175181e-09, 6.013818e-08, -3.07158e-08, 3.974361e-08, 1.740335e-08, 
    -1.186947e-09, -7.425683e-09, 2.040076e-08, -2.216939e-08, 1.2339e-09, 
    -1.860542e-08, -2.297577e-09, 1.291752e-09, -2.053162e-08, 5.98741e-09, 
    2.468122e-08, -3.069374e-09, 1.539402e-08, 1.703221e-09, -1.57429e-08, 
    -2.513525e-08, 5.35664e-08, 6.266177e-09, -9.37281e-09, -9.539498e-10, 
    4.634543e-09, -9.211362e-09, 1.485675e-08, -1.061051e-09, -3.017008e-09, 
    5.50159e-10, 7.760178e-08, 1.017719e-08, 1.53774e-08, -9.261022e-09, 
    -3.290609e-09, 5.969468e-09, -5.305196e-10, -2.1473e-08, 8.706366e-10, 
    -1.359234e-08, 1.021743e-08, 2.827562e-08, 1.516935e-08, 8.759173e-09, 
    -2.191769e-09, 2.356222e-08, -3.70116e-08, -1.899707e-10, 2.231648e-08, 
    2.330012e-10, 2.283116e-10, -2.703547e-08, 4.727556e-09, 2.928766e-08, 
    -1.740136e-08, -2.061678e-08, -1.173362e-09, 7.607923e-10, -2.864908e-10, 
    4.790991e-09, -5.415473e-10, -1.749811e-09, -9.261354e-09, -1.726497e-08, 
    5.17889e-09, 4.448966e-08, -5.550319e-09, 1.138617e-08, 9.741768e-09, 
    2.426891e-08, -1.630065e-09, -3.292945e-08, -3.814648e-09, -3.503192e-09, 
    -1.522778e-09, 1.238319e-08, 7.944934e-11, -7.949943e-10, 1.699254e-08, 
    3.343018e-09, -2.769241e-09, -1.107395e-08, 1.300782e-08, 7.594679e-09, 
    3.134232e-09, -6.575135e-09, 5.379718e-09, 1.21554e-09, -7.053018e-09, 
    -7.374751e-10, 1.218019e-09, 3.676526e-10, 3.602452e-12, -3.613309e-09,
  2.922889e-09, -1.621117e-09, -4.521155e-09, -1.318256e-09, 2.063416e-10, 
    -2.30898e-10, 6.950074e-09, -3.872685e-09, 9.592441e-09, 7.287326e-10, 
    3.731202e-10, -4.756089e-10, -5.688548e-09, -1.072624e-08, 2.927612e-08, 
    -3.247226e-09, -8.871444e-09, 1.457352e-09, 5.365308e-09, 8.429424e-09, 
    3.364164e-09, -1.67359e-08, -1.483613e-09, 9.609323e-09, 6.233449e-10, 
    1.161027e-09, 6.73345e-08, -8.125312e-09, -3.983911e-08, 1.863714e-08, 
    -2.83984e-09, -3.000764e-09, 3.864756e-08, -4.057688e-08, 2.193701e-09, 
    -2.619885e-08, -3.516971e-09, 1.873644e-09, -1.231041e-08, 1.519703e-08, 
    3.359542e-08, 6.792391e-09, 1.925926e-08, 2.115081e-09, -2.640155e-08, 
    -1.28457e-08, 4.924973e-08, 1.081439e-08, -1.787624e-08, -1.487457e-09, 
    1.259713e-08, -1.118207e-08, 2.555255e-08, -2.815807e-09, -3.158701e-09, 
    5.359198e-10, 1.321551e-07, 1.47243e-08, 2.750543e-08, -1.534868e-08, 
    -7.085248e-09, 4.802416e-09, 3.438174e-09, -2.506317e-08, -1.510898e-10, 
    -4.220311e-08, 6.915116e-09, 1.591388e-08, 2.057965e-08, 7.485653e-09, 
    -3.976879e-09, 2.350703e-09, -4.875562e-08, 2.121226e-09, 3.613708e-08, 
    1.652438e-10, 3.712017e-10, -3.265455e-08, 5.051401e-09, 3.434496e-08, 
    -1.725834e-08, -1.424563e-08, -2.898446e-09, 1.317119e-09, -4.261494e-09, 
    3.752632e-09, 8.528218e-10, -5.099423e-10, -1.347025e-08, -1.957201e-08, 
    1.341903e-09, 6.93906e-08, -3.972787e-09, 6.57256e-08, 9.760299e-09, 
    3.196906e-08, -1.346848e-09, -9.272469e-09, -5.065772e-09, -4.971343e-09, 
    -2.557613e-09, 5.145761e-09, -6.316192e-10, 4.888001e-10, 9.254904e-09, 
    -8.03027e-10, -7.324104e-09, 9.886321e-09, 2.254251e-08, 5.173717e-09, 
    6.771188e-10, -4.938556e-09, 3.514174e-09, -3.299192e-10, -1.541991e-08, 
    -1.141819e-09, 1.804707e-09, 4.761027e-10, 4.337863e-11, -2.980755e-09,
  2.579952e-09, -1.979743e-09, -7.14067e-10, -1.144542e-08, 1.141302e-09, 
    1.226397e-09, 6.966445e-09, -2.106788e-08, 4.285084e-09, -2.85371e-09, 
    -4.938556e-10, 6.858727e-10, -1.950752e-09, -4.460901e-09, -1.233445e-08, 
    -2.111939e-09, -1.117693e-08, 4.259618e-09, 6.38989e-09, 1.158804e-08, 
    1.089933e-08, -2.778449e-09, -6.9561e-09, 1.377481e-08, -1.301714e-11, 
    6.488108e-10, 4.516761e-08, 1.75616e-08, -3.476578e-08, 1.389498e-08, 
    -2.870593e-09, -3.205685e-09, 6.673412e-08, -8.187226e-08, 9.238931e-09, 
    -3.786772e-08, -5.942769e-09, 2.447102e-09, 1.432494e-08, 2.078806e-08, 
    3.863926e-08, 5.185086e-09, 1.936232e-08, 1.472817e-09, -2.120782e-08, 
    1.277607e-08, 4.225126e-08, 1.203895e-08, -1.145866e-08, -2.293046e-09, 
    1.841965e-08, -7.054325e-09, 4.011441e-08, -1.445449e-09, -9.616141e-09, 
    3.854836e-10, 1.549641e-07, 1.119551e-08, 3.255179e-08, -2.228014e-08, 
    3.189484e-10, 6.383686e-09, 6.43621e-09, -3.116362e-08, -4.771743e-09, 
    -8.677438e-08, 8.713528e-09, -4.446974e-09, 3.111461e-08, -1.288896e-08, 
    -1.417163e-09, -2.859662e-08, -5.119722e-08, -2.681361e-09, 4.341353e-08, 
    -2.513048e-10, 9.964793e-10, -3.746263e-08, 3.23225e-09, 1.63152e-08, 
    -1.484028e-08, 6.285123e-09, -4.729657e-09, 2.031356e-09, -2.537774e-09, 
    -1.421711e-09, 8.699885e-10, 3.27384e-09, -1.525821e-08, -2.052167e-08, 
    -2.668742e-09, 9.619698e-08, -2.069811e-10, 1.510424e-07, 9.628309e-09, 
    3.975641e-08, -1.777016e-09, 3.1399e-08, -5.15746e-09, -5.913717e-09, 
    -3.118828e-09, -1.045883e-09, -1.23093e-09, 1.167411e-09, 3.594891e-09, 
    -2.812044e-10, -2.487752e-09, 1.160419e-08, 1.402196e-08, 1.599972e-09, 
    -2.382194e-09, -1.130729e-09, 6.674554e-10, -8.110987e-10, -2.501775e-08, 
    -1.480089e-09, 2.322544e-09, 6.403944e-10, 6.948753e-11, -5.672405e-10,
  5.286438e-11, -1.638682e-09, 1.58758e-08, -3.747857e-08, -3.752803e-10, 
    -4.930598e-10, 6.511982e-10, -2.64381e-08, -4.35989e-10, -7.722974e-09, 
    -5.693437e-10, 4.136609e-09, 4.561116e-10, 3.522814e-09, -1.322019e-08, 
    -1.993815e-09, -1.312008e-08, 8.820507e-09, 7.776507e-09, 1.076887e-08, 
    3.647676e-08, 4.615345e-09, -1.411217e-08, 7.960125e-09, -1.961098e-10, 
    -2.373781e-10, -9.703058e-09, 3.045704e-08, 1.588886e-07, 9.743417e-09, 
    7.604865e-08, -8.170105e-09, 5.502523e-08, -1.126059e-07, 1.61973e-08, 
    -4.870333e-08, -7.258472e-09, 3.018755e-09, -5.325774e-09, 2.201029e-08, 
    3.292741e-08, 5.925699e-09, 1.633475e-08, -4.49079e-10, -1.490207e-08, 
    9.152927e-09, 4.142396e-08, 3.4219e-08, 2.157201e-08, -3.360384e-09, 
    2.123876e-08, -1.047272e-08, 6.274748e-08, -3.465812e-09, -1.063321e-08, 
    6.423306e-11, 1.537857e-07, 6.541439e-09, 3.125019e-08, -2.228785e-08, 
    2.061438e-08, 9.004452e-09, 5.300762e-09, -4.094586e-08, -7.91299e-09, 
    -5.984521e-08, 1.15976e-07, -2.718741e-08, 3.521927e-08, -5.705465e-08, 
    -5.178094e-09, -5.467859e-08, -3.340915e-08, -8.119741e-09, 4.036431e-08, 
    -8.735697e-10, 9.372059e-10, -4.010622e-08, -4.888562e-10, 1.330591e-09, 
    -1.193229e-08, 3.126856e-08, -6.314167e-09, 1.435751e-09, -4.552589e-09, 
    -1.796025e-08, 4.120125e-09, 6.665459e-09, -6.372566e-09, -2.906035e-08, 
    -8.998086e-09, 1.11353e-07, 1.823423e-09, 1.981091e-07, 3.349442e-09, 
    4.418859e-08, 3.445166e-09, 6.215635e-08, -4.070671e-09, -6.367509e-09, 
    -2.603542e-09, -4.033751e-10, -1.385104e-09, 1.860165e-09, -3.843297e-09, 
    7.423751e-10, -5.764718e-09, -1.443993e-08, 5.257903e-09, -1.414946e-09, 
    -6.381356e-09, 8.119514e-10, -1.091848e-09, -1.723265e-09, -1.747958e-08, 
    -1.763283e-09, 2.82671e-09, 8.480399e-10, 3.177547e-11, 2.065349e-09,
  1.575188e-08, 1.349804e-09, 4.9449e-08, -7.163351e-08, -8.770598e-09, 
    -7.396579e-09, -1.50294e-10, -1.18041e-08, -1.800333e-08, -7.609628e-09, 
    1.358671e-09, 5.513812e-09, 1.005787e-09, 2.249681e-08, -5.456968e-11, 
    -3.034256e-09, -1.653036e-08, 4.505011e-09, 3.267601e-09, 5.400807e-09, 
    4.476749e-08, -1.133503e-08, 1.648232e-09, -2.043635e-09, 1.301714e-09, 
    -3.438231e-09, 1.659828e-10, 3.356433e-08, 1.712463e-07, 1.089222e-08, 
    4.368235e-08, -2.23838e-08, 6.921391e-08, -6.578364e-08, 1.620197e-08, 
    -4.809522e-08, -6.421124e-09, 4.462848e-09, -3.338425e-08, 3.52821e-08, 
    1.598464e-08, 7.974336e-09, 1.844131e-08, -1.366271e-09, -1.155774e-08, 
    -3.117293e-09, 4.413175e-08, 7.454676e-08, 3.762634e-08, -4.605198e-09, 
    2.228552e-08, -2.927459e-08, 1.020936e-07, -8.895291e-09, -8.108873e-09, 
    -4.614549e-10, 1.164492e-07, 1.226036e-08, 3.714302e-08, -1.247041e-08, 
    1.511319e-08, 5.807237e-09, 2.384581e-09, -5.259303e-08, -1.603962e-08, 
    -4.328388e-08, 1.173606e-07, -4.862079e-08, 3.304035e-08, -3.728564e-08, 
    -1.204637e-08, -9.797054e-08, -1.574369e-08, -5.27541e-09, 4.414314e-08, 
    -1.966214e-09, 5.108944e-10, -3.701115e-08, -3.679483e-09, -1.139028e-09, 
    -9.44766e-09, 3.651442e-08, -7.934375e-09, -1.070589e-09, 1.258172e-09, 
    3.734272e-08, 1.350395e-08, 5.366815e-09, -8.068863e-09, -4.306293e-08, 
    -9.755354e-09, 1.207995e-07, 1.945494e-09, 1.898775e-07, -1.044521e-08, 
    4.356691e-08, 1.917972e-08, 2.863328e-08, -3.041919e-09, -7.893595e-09, 
    6.034497e-10, -9.61947e-10, -6.458386e-09, 1.046416e-10, 2.477918e-09, 
    2.089041e-08, -1.614342e-08, -3.34627e-08, -3.583523e-09, -3.411969e-09, 
    -9.461701e-09, 5.915126e-10, -1.230546e-09, -2.809884e-09, 1.085255e-09, 
    -2.139779e-09, 3.335728e-09, 5.149907e-10, -2.98499e-11, 4.70834e-09,
  8.436774e-08, 2.908507e-09, 6.480906e-08, -7.159446e-08, -2.766507e-08, 
    -6.146877e-09, 2.486274e-09, 1.519936e-09, -2.333996e-08, 6.195933e-12, 
    3.981938e-09, 4.327205e-09, 2.285276e-09, 3.776319e-08, 2.094396e-09, 
    -5.078959e-09, -2.335487e-08, 2.59314e-09, -1.455018e-08, -2.110426e-09, 
    3.712159e-09, -2.464623e-08, -2.583971e-08, -3.338243e-09, -8.95551e-09, 
    -7.714505e-09, 6.629648e-10, 2.89869e-08, 9.757667e-08, 1.288021e-08, 
    2.356234e-08, -9.285856e-08, 8.037415e-08, 3.386521e-08, 7.170058e-09, 
    -3.702695e-08, -2.463833e-09, 6.861356e-09, -4.195442e-09, 2.623142e-08, 
    -7.362019e-10, 7.234064e-09, 1.830793e-08, 8.70374e-10, -2.999457e-09, 
    -1.769621e-08, 4.722705e-08, 1.037611e-07, 4.633404e-08, -5.896013e-09, 
    2.118523e-08, -5.388057e-08, 1.740573e-07, -1.231614e-08, 2.762693e-09, 
    -1.231854e-09, 1.046263e-07, 2.814284e-08, 5.052566e-08, 7.69748e-09, 
    2.391573e-09, 2.103036e-09, -1.151079e-10, -7.013981e-08, -2.858727e-08, 
    -3.846748e-08, 1.478313e-07, -5.951648e-08, 2.830558e-08, 4.218651e-08, 
    8.694713e-09, -1.037359e-07, -1.846621e-08, -3.908042e-09, 6.98971e-08, 
    -2.964669e-09, 7.499068e-10, -3.152968e-08, -5.594987e-09, 9.985075e-08, 
    -6.356402e-09, 1.494062e-08, -9.027758e-09, -5.199297e-09, 7.971551e-09, 
    1.673487e-08, -5.499317e-09, 4.31811e-09, -1.673325e-08, -5.071882e-08, 
    -6.273524e-09, 1.228576e-07, 1.744866e-09, 1.509177e-07, -8.223043e-08, 
    3.788982e-08, 5.707133e-08, 2.324322e-08, -1.141814e-09, -1.2716e-08, 
    1.828596e-09, -5.732595e-09, 4.239055e-09, -4.280679e-09, 4.067766e-08, 
    5.202418e-08, -2.245434e-08, -5.260819e-08, -9.821349e-09, 9.771384e-11, 
    -7.871392e-09, -1.19195e-09, -8.519123e-10, -2.400554e-09, 5.211575e-09, 
    -2.574836e-09, 3.444129e-09, 3.021654e-10, -1.069296e-10, -5.416553e-09,
  9.437508e-08, 6.895107e-10, 6.025982e-08, 4.192384e-08, -3.163109e-08, 
    -3.858645e-09, 4.530989e-09, 1.711589e-08, -1.115575e-08, 4.452659e-09, 
    3.999503e-09, 3.040668e-09, 1.610715e-09, 5.039772e-08, 1.825128e-09, 
    -7.598139e-09, -3.05052e-08, 1.494601e-08, -3.210945e-08, 2.599904e-09, 
    -2.287572e-08, -1.118406e-08, -3.311129e-08, -5.292839e-08, -2.05257e-08, 
    -1.300805e-09, 4.733977e-08, 3.31363e-09, 4.537821e-08, 2.337504e-08, 
    2.491618e-08, -3.948844e-08, 1.652052e-08, -7.172844e-09, -1.458216e-08, 
    -2.723345e-08, 4.018716e-09, 1.024809e-08, 1.886383e-08, 1.833359e-08, 
    -2.612637e-08, 3.714035e-09, 1.067917e-08, 5.718164e-10, -1.083754e-08, 
    -4.58158e-08, 5.034479e-08, 9.400685e-08, 5.029138e-08, -7.006932e-09, 
    1.883723e-08, -6.253993e-08, 2.494016e-07, -1.154415e-08, 1.739705e-08, 
    -8.857342e-10, 1.000932e-07, 3.064604e-08, 4.518934e-08, 3.34086e-08, 
    1.728495e-09, 4.088179e-10, 1.520334e-09, -8.871314e-08, -4.863864e-08, 
    -3.84432e-08, 1.212168e-07, -5.343873e-08, 2.381955e-08, 6.796381e-08, 
    1.216893e-08, -1.348969e-07, -3.657556e-08, -6.766982e-09, 8.40198e-08, 
    -1.074682e-09, 1.522537e-09, -1.803764e-08, -7.434733e-09, -2.973547e-08, 
    -6.344806e-09, -5.356148e-09, -1.083231e-08, -5.382617e-09, 3.632863e-09, 
    2.432432e-08, -9.52241e-10, 1.678586e-09, -1.5541e-08, -5.286455e-08, 
    -1.717694e-09, 1.126154e-07, 2.243866e-09, 1.219779e-07, -6.812922e-08, 
    2.574443e-08, 8.422287e-08, 5.414768e-08, 1.205876e-09, -1.970509e-08, 
    4.231765e-09, -6.277254e-09, 5.023537e-10, -1.472211e-08, 6.735297e-08, 
    5.526886e-08, -2.883235e-08, -6.07821e-08, -2.010177e-08, 3.83352e-10, 
    -3.818286e-09, -2.263505e-09, -3.284072e-09, -3.17641e-10, -1.538751e-09, 
    -2.770378e-09, 3.296819e-09, -4.000604e-10, -1.874625e-10, -1.836258e-08,
  3.132891e-08, -2.189495e-09, 4.196454e-08, 1.361424e-07, -1.138892e-08, 
    1.003855e-10, 1.284309e-08, 1.116427e-08, 1.912667e-08, 3.320565e-09, 
    4.763479e-10, -2.921752e-11, 1.694957e-09, 4.342974e-08, -2.306365e-09, 
    -1.639575e-08, -4.318165e-08, 3.426288e-08, -1.10247e-07, 2.168929e-08, 
    -3.790171e-08, 6.031428e-09, 1.07691e-08, -1.513524e-08, 2.934485e-09, 
    4.803042e-09, 9.092753e-08, -1.001695e-09, 3.327193e-08, 3.62669e-08, 
    4.842911e-08, 7.127528e-08, 5.384209e-09, -8.887071e-08, -4.054198e-08, 
    -3.020955e-08, 1.017087e-08, 1.506548e-08, 5.597178e-08, -5.865161e-09, 
    -6.476441e-08, 1.693934e-11, 5.993286e-09, -3.498e-09, -3.256105e-08, 
    -8.919346e-08, 6.415331e-08, 3.446866e-08, 5.19349e-08, -6.881464e-09, 
    1.468432e-08, -4.617345e-08, 2.978981e-07, -7.568474e-09, 4.240254e-08, 
    -5.853735e-10, 9.777375e-08, 2.552758e-08, 3.293868e-08, 3.990117e-08, 
    9.466703e-10, 2.455636e-11, -6.161486e-09, -9.602773e-08, -6.859646e-08, 
    -6.898847e-08, 1.046782e-07, -4.762126e-08, 1.684532e-08, 8.668894e-08, 
    9.798327e-09, -1.739028e-07, -4.687797e-08, -1.775038e-08, 6.173186e-08, 
    -7.491963e-11, 3.63903e-09, 4.514646e-09, -9.139776e-09, -1.32977e-07, 
    -7.764697e-09, -1.456689e-09, -2.161516e-08, -4.705043e-09, -5.20015e-09, 
    -5.814525e-08, 1.038757e-09, -1.244757e-09, -8.068772e-09, -5.069165e-08, 
    -1.885496e-09, 7.470107e-08, 2.562217e-09, 1.051824e-07, -9.010478e-09, 
    1.138999e-08, -8.890401e-09, 5.10471e-08, -1.052967e-09, -2.609513e-08, 
    -1.280262e-08, 4.258482e-09, -8.914391e-09, -2.384543e-08, 7.740368e-08, 
    3.048706e-08, -2.459433e-08, -5.77802e-08, -2.440561e-08, -4.314188e-09, 
    7.762878e-09, -4.501999e-10, -3.490413e-09, -1.455192e-11, -2.39163e-09, 
    -2.755246e-09, 3.339323e-09, -8.192522e-10, -2.731113e-10, -7.298695e-09,
  -6.582241e-08, -1.581839e-09, 1.609612e-08, 1.123287e-07, -1.518345e-08, 
    1.000819e-08, 2.165643e-08, 1.776584e-09, 2.862953e-08, 4.912977e-09, 
    1.815579e-10, -6.551772e-10, 9.791961e-09, 7.507879e-10, -7.379526e-09, 
    -2.637495e-08, -4.324139e-08, 5.985504e-08, -2.158056e-07, 3.165769e-08, 
    -3.799676e-08, 5.22266e-09, 3.178434e-08, 2.484342e-08, 1.485807e-08, 
    2.034312e-09, 4.385345e-08, 2.298475e-08, 3.531397e-08, 3.897878e-08, 
    2.647118e-08, 5.300058e-08, 2.189518e-08, -7.147071e-08, -6.250525e-08, 
    -2.774038e-08, 1.362613e-08, 2.022597e-08, 8.526058e-08, -5.153927e-08, 
    -1.315289e-07, 3.200057e-09, 4.576407e-09, -7.265617e-09, -3.165849e-08, 
    -1.110869e-07, 1.173366e-07, -4.459207e-08, 5.182562e-08, -5.925934e-09, 
    1.013052e-08, -3.424805e-08, 3.053579e-07, -7.795075e-09, 6.576435e-08, 
    -1.149374e-09, 9.893256e-08, 9.234339e-09, 4.231033e-08, 3.226633e-08, 
    -1.647095e-09, -3.956302e-11, 1.063245e-08, -8.136408e-08, -7.668962e-08, 
    -1.148549e-07, 3.701575e-08, -3.080459e-08, 1.135277e-08, 6.960818e-08, 
    8.313737e-08, -1.649574e-07, -4.950698e-08, -1.723834e-08, 5.111901e-08, 
    -8.352458e-09, 5.343296e-09, 4.362704e-08, -1.025126e-08, -3.421894e-08, 
    -1.007277e-08, -5.548884e-10, -4.402688e-08, -2.502247e-09, 
    -7.631002e-09, 2.642321e-08, -1.054807e-07, 3.232799e-09, 3.150383e-09, 
    -4.224194e-08, 1.150511e-10, 2.770321e-08, 1.758593e-09, 1.223538e-07, 
    -1.180933e-08, -8.780852e-09, -2.15161e-08, 7.738208e-09, -4.593517e-09, 
    -3.175071e-08, -3.511195e-08, 1.003482e-08, -4.487198e-09, -3.113963e-08, 
    3.856871e-08, 1.180865e-09, -2.166053e-08, -4.028755e-08, -1.842898e-08, 
    -1.287708e-08, 1.117326e-08, 3.799414e-10, -4.452431e-09, -6.751293e-09, 
    2.481784e-10, -2.612956e-09, 3.762224e-09, -1.006029e-09, -3.886811e-10, 
    -2.465868e-10,
  -5.06314e-08, -4.455956e-10, 3.76366e-09, 2.463361e-08, -1.659822e-08, 
    1.652353e-08, 3.421945e-08, -2.104372e-08, 2.037211e-09, -3.723528e-09, 
    -3.049024e-09, 3.105356e-10, 1.937514e-08, -3.308952e-08, -9.585563e-09, 
    -3.395159e-08, -4.632575e-08, 8.231353e-08, -2.48403e-07, 3.652525e-08, 
    -3.782606e-08, 1.765727e-09, 1.410996e-08, 9.252005e-09, 5.29252e-09, 
    -8.985751e-09, 2.883218e-08, 3.032034e-08, 2.637518e-08, 3.917881e-08, 
    4.741383e-08, 2.235316e-08, 4.484394e-08, 4.391831e-08, -8.778505e-08, 
    -2.228245e-08, 1.450824e-08, 2.437632e-08, 9.654929e-08, -5.9751e-08, 
    -1.979858e-07, 6.278754e-09, 4.973316e-09, -9.641804e-09, -3.17213e-08, 
    -1.108745e-07, 1.435089e-07, -1.260082e-07, 3.766414e-08, -5.967323e-09, 
    7.976041e-09, -3.034705e-08, 2.569309e-07, -9.760913e-09, 8.422347e-08, 
    -1.335593e-09, 1.057521e-07, -2.792671e-09, 6.378022e-08, 2.507043e-08, 
    -1.416595e-09, -3.099382e-08, 1.141775e-07, -7.10288e-08, -6.217395e-08, 
    -1.284132e-07, -2.005635e-08, -4.822027e-10, 7.211895e-09, 6.024874e-08, 
    -9.08214e-08, -1.607368e-07, -3.630174e-08, -5.133529e-10, 7.875237e-08, 
    -2.203461e-08, 4.448239e-09, 7.014958e-08, -1.153809e-08, 4.923606e-09, 
    -1.171924e-08, -2.659002e-08, -5.649315e-08, -2.979675e-09, 
    -1.158867e-09, 6.20542e-08, -1.502283e-07, 1.005827e-08, -1.791427e-08, 
    -2.879688e-08, 1.840743e-08, 4.395827e-09, -1.349434e-09, 1.261918e-07, 
    -2.168605e-08, -2.470813e-08, 2.509561e-08, -1.937343e-08, -2.211863e-08, 
    -3.699805e-08, 4.187149e-08, -2.18121e-09, -1.538659e-09, -2.907866e-08, 
    1.705774e-08, 7.043525e-09, -3.526583e-08, -2.306132e-08, -8.661516e-09, 
    -6.667449e-09, 3.660659e-09, -2.612012e-09, -1.055884e-08, -2.174767e-08, 
    1.256751e-09, -2.167235e-09, 6.565401e-09, -1.14148e-09, -5.276988e-10, 
    -7.747298e-08,
  -4.434037e-08, 6.998562e-10, 2.966999e-09, -2.055629e-08, 1.850935e-09, 
    1.348644e-08, 5.343918e-08, -3.607488e-08, -2.740353e-08, -6.845198e-09, 
    -1.481567e-09, -9.081305e-10, 1.349008e-08, -3.768127e-08, -8.372695e-09, 
    -3.282339e-08, -5.487212e-08, 7.560988e-08, -1.532486e-07, 1.586523e-08, 
    -3.222772e-08, 2.524712e-08, 1.188596e-09, -2.915499e-09, -2.190518e-09, 
    -4.882725e-08, 1.246474e-08, 2.438344e-08, 8.737175e-09, 3.958792e-08, 
    5.579818e-08, 8.26401e-09, 4.899448e-08, 9.451048e-08, -1.272291e-07, 
    -1.673243e-08, 2.741206e-09, 2.785005e-08, 1.083662e-07, 1.578925e-08, 
    -1.144097e-07, 4.301228e-09, 2.493721e-09, -1.017125e-08, -2.866796e-08, 
    -9.620942e-08, 1.581632e-07, -1.455242e-07, -9.041514e-09, -8.129355e-09, 
    7.627506e-09, -3.105038e-08, 1.835857e-07, -1.05684e-08, 9.894738e-08, 
    -1.065587e-09, 1.123458e-07, -6.697597e-08, 8.317552e-08, 2.19827e-08, 
    1.012836e-09, -5.95262e-08, 1.190301e-08, -7.727235e-08, -4.806334e-08, 
    -1.090341e-07, 3.567402e-08, 1.380192e-08, 1.964054e-09, 7.19599e-08, 
    4.222954e-08, -1.171428e-07, -4.861874e-08, 2.547722e-10, 1.052443e-07, 
    -3.409332e-08, 3.343388e-09, 8.822627e-08, -1.017719e-08, -1.281103e-08, 
    -1.279153e-08, -1.053678e-07, -3.46642e-08, -6.310756e-09, -2.924253e-09, 
    5.769698e-08, -1.625472e-08, 2.881814e-08, -5.737693e-08, -3.392984e-08, 
    1.461319e-08, -3.196455e-08, -3.329689e-09, 1.206137e-07, -4.365643e-08, 
    -2.89527e-08, -1.024284e-08, 1.432966e-08, -3.146772e-08, -3.948819e-08, 
    6.29027e-08, -3.087788e-08, 1.386979e-11, -1.821871e-08, 4.703418e-08, 
    3.905188e-08, -1.973274e-08, -2.686386e-08, 7.391009e-09, 2.190711e-08, 
    -1.764533e-09, -5.086349e-09, -1.657907e-08, -3.916591e-08, 
    -3.808395e-09, -1.682508e-09, 1.117094e-08, -1.219234e-09, -6.703615e-10, 
    -8.786822e-08,
  -4.118613e-08, 2.170054e-09, 3.514515e-09, -1.882358e-08, 1.749618e-08, 
    2.100558e-08, 6.71514e-08, -2.173533e-08, -4.609285e-08, -1.898445e-08, 
    3.364676e-09, -5.950369e-10, -2.031686e-08, 1.141223e-08, 3.648211e-09, 
    -3.647798e-08, -6.013394e-08, 4.728452e-08, -6.654082e-08, -5.147763e-08, 
    -1.684953e-09, 1.052703e-07, -1.711783e-09, -9.063115e-10, -3.918308e-08, 
    -1.752934e-07, 1.340118e-08, 1.641331e-08, 2.232355e-09, 3.646085e-08, 
    5.657216e-08, 9.48819e-09, 3.692719e-08, 9.569442e-08, -1.344516e-07, 
    -3.631249e-08, -3.843638e-10, 3.062878e-08, 1.178768e-07, 7.419648e-08, 
    -7.975984e-08, 1.444164e-09, 2.297696e-09, -7.554883e-09, -2.474269e-08, 
    -1.11192e-07, 1.607551e-07, -5.155698e-08, -5.860647e-08, -1.019166e-08, 
    7.411927e-09, -4.123751e-08, 1.109936e-07, -1.100382e-08, 1.037172e-07, 
    -5.375114e-10, 1.032494e-07, -6.889738e-08, 9.591957e-08, -5.250655e-09, 
    2.49986e-09, -3.693469e-08, 7.173878e-08, -9.088217e-08, -6.181026e-08, 
    -8.669667e-08, -2.147158e-08, 3.090656e-08, 3.931291e-10, 6.969128e-08, 
    1.389333e-07, -5.812865e-08, -1.018235e-07, -9.645532e-09, 1.076045e-07, 
    -3.934213e-08, 7.906294e-09, 8.203779e-08, -1.42343e-09, -5.491279e-08, 
    -1.181905e-08, -1.613362e-07, 1.073715e-08, -1.087803e-07, -5.182983e-08, 
    4.006506e-08, 1.263905e-07, 5.773313e-08, -6.496914e-08, -4.05833e-08, 
    8.013217e-09, -9.039386e-08, -4.661757e-09, 1.130092e-07, -8.831796e-08, 
    1.236755e-07, -7.863476e-08, 1.115893e-08, -4.246465e-08, -3.755115e-08, 
    -1.476972e-07, -4.298303e-08, -2.723354e-09, -8.088612e-09, -2.56822e-08, 
    4.00729e-08, -1.885473e-08, -2.796378e-08, 1.947683e-08, 3.669845e-08, 
    -5.623747e-09, -3.467107e-09, -1.652688e-08, -4.919946e-08, 
    -6.895561e-09, -9.258088e-10, 1.614173e-08, -1.051642e-09, -7.717347e-10, 
    -7.344909e-08,
  -4.035587e-08, 6.87362e-09, 4.821572e-09, 1.114165e-08, 4.048684e-08, 
    2.778495e-08, 7.951121e-08, 3.193691e-09, -2.813761e-08, -3.733851e-08, 
    1.392209e-09, -2.194304e-08, -2.500849e-08, -2.808417e-08, -8.960797e-10, 
    -3.376692e-08, -5.10953e-08, 5.230788e-08, -6.720835e-08, -1.406823e-07, 
    5.902348e-08, 7.919311e-08, -9.420887e-09, -1.391413e-09, -7.068491e-08, 
    -1.457366e-07, 3.076252e-08, 1.502758e-08, -1.270678e-09, 3.672653e-08, 
    7.891822e-08, 1.221713e-08, 2.304466e-08, 3.560228e-08, -1.259697e-07, 
    -3.663604e-08, -1.274159e-08, 3.256538e-08, 1.201781e-07, 1.11299e-07, 
    -1.049233e-07, -4.409571e-09, 1.496468e-08, 2.927115e-09, -1.60361e-08, 
    -1.382102e-07, 9.759168e-08, 6.614835e-08, -8.391628e-08, -1.10848e-08, 
    6.600914e-09, -2.340323e-08, 5.599843e-08, -8.893084e-09, 9.82738e-08, 
    -4.025708e-09, 9.640587e-08, 3.164455e-08, 1.04542e-07, -4.693335e-08, 
    1.802277e-09, -2.066668e-08, 3.924083e-08, -1.081005e-07, -2.291047e-08, 
    -4.348271e-08, -6.48015e-11, 2.666854e-08, -1.70553e-09, 6.13835e-08, 
    1.550815e-07, -1.901298e-07, -6.93035e-08, -8.602342e-09, 9.198033e-08, 
    -3.181515e-08, 7.573973e-09, 8.198774e-08, 1.020572e-08, 4.409799e-09, 
    -7.569497e-09, -1.944431e-07, 4.170596e-08, -1.407017e-07, -2.433353e-08, 
    1.824894e-07, 5.608308e-08, 8.187169e-08, -4.72311e-08, -3.182532e-08, 
    7.124413e-09, -1.156722e-07, -5.227605e-09, 8.913392e-08, -1.001603e-07, 
    9.991372e-08, -1.34354e-07, -2.091588e-08, -5.488369e-08, -3.001069e-08, 
    -3.142679e-08, -3.250548e-08, -2.526292e-09, -4.902304e-09, 
    -2.259321e-08, -2.060085e-08, -1.980254e-08, -1.123567e-09, 1.840408e-08, 
    2.897968e-08, -2.3501e-08, -2.589331e-09, -7.112249e-09, -5.49868e-08, 
    -5.054972e-09, -9.056066e-10, 1.849791e-08, -7.123582e-10, -8.995826e-10, 
    -9.718713e-08,
  -2.000615e-08, 1.620401e-08, 5.903644e-09, 4.738604e-08, 7.246604e-08, 
    3.227342e-08, 8.824907e-08, 2.564548e-08, 1.004764e-09, -2.510671e-08, 
    -9.406676e-09, -6.261632e-08, 2.148113e-09, -5.327934e-08, 6.756295e-09, 
    -4.460431e-08, -3.586068e-08, 4.625997e-08, -5.100489e-08, -1.924548e-08, 
    1.105263e-07, -4.988794e-08, -9.653797e-08, -4.985918e-08, -5.183142e-08, 
    -1.198105e-07, 3.233151e-08, 1.414242e-08, -9.486712e-09, 4.713854e-08, 
    9.412759e-08, 6.802452e-09, 1.563819e-08, -4.420951e-08, -1.119666e-07, 
    -2.832508e-08, -2.058893e-08, 3.279297e-08, 1.138021e-07, 1.262397e-07, 
    -1.290268e-07, -2.313785e-07, -6.984536e-08, 2.27065e-08, -3.171499e-08, 
    -1.101622e-07, 8.000188e-08, 1.405139e-07, -7.451247e-08, -9.228515e-09, 
    5.741967e-09, -1.086055e-07, 2.304156e-08, -1.5003e-08, 7.647814e-08, 
    -7.573078e-09, 8.540906e-08, 1.001346e-07, 1.072069e-07, -6.793354e-08, 
    -9.112e-10, -4.192611e-08, 2.993204e-08, -1.136794e-07, -3.476408e-09, 
    -2.140996e-08, 6.900564e-09, 2.07491e-08, 1.126068e-09, 4.739115e-08, 
    6.110577e-08, -1.994059e-07, -2.054935e-08, -1.096237e-08, 6.384157e-08, 
    -2.445279e-08, -4.619778e-09, 7.45068e-08, 2.294744e-08, -2.052218e-08, 
    2.071147e-09, -1.892835e-07, 6.278356e-08, -1.091333e-07, 1.034927e-07, 
    2.582193e-07, -5.052516e-08, 7.607866e-08, -3.719134e-08, -2.289215e-08, 
    -5.657739e-09, -1.089868e-07, -4.660336e-09, 2.626103e-08, -8.35613e-08, 
    7.902747e-08, -1.711474e-07, -2.978709e-08, -6.365724e-08, -3.311172e-08, 
    1.027831e-08, -1.885129e-08, -1.054644e-09, -1.045429e-09, 7.393828e-08, 
    -4.406911e-08, -1.982926e-08, 3.602031e-08, 8.017537e-09, 1.236572e-08, 
    -6.458845e-08, -2.941988e-09, 2.66823e-10, -4.736069e-08, -1.310696e-09, 
    4.186859e-10, 1.371951e-08, -8.001528e-10, -1.030251e-09, -1.622575e-07,
  -3.555272e-09, 3.174415e-08, 3.87405e-09, 3.251233e-08, 4.055715e-08, 
    3.558631e-08, 8.981471e-08, 3.402334e-08, 2.168605e-08, -5.158711e-09, 
    -5.914893e-08, -4.696557e-08, 3.865358e-08, -2.878954e-08, 1.142433e-08, 
    -3.796242e-08, -1.883368e-08, 7.95701e-08, -5.788124e-08, -2.343853e-08, 
    1.194152e-07, -1.677626e-08, -1.433071e-07, -1.409256e-07, 1.596987e-08, 
    -9.056947e-08, 4.777752e-08, 1.340999e-08, -1.73273e-08, 8.690591e-08, 
    8.085857e-08, 6.521816e-09, 1.585937e-08, -1.295182e-07, -1.17262e-07, 
    -2.879682e-08, -2.701148e-08, 3.183513e-08, 9.629235e-08, 1.524607e-07, 
    -1.034492e-07, -1.579156e-07, -2.052816e-07, 4.713799e-08, -2.112228e-08, 
    -7.558214e-08, 1.628479e-08, 2.059143e-07, -5.587768e-08, -6.235396e-09, 
    5.43524e-09, -1.893886e-07, 5.009644e-09, -1.071754e-08, 4.321952e-08, 
    -4.28588e-09, 6.797808e-08, 1.519774e-07, 1.106053e-07, -8.146137e-08, 
    -2.238096e-09, -8.75919e-08, 4.128134e-08, -1.248407e-07, 2.246487e-08, 
    -3.180247e-08, 2.42739e-08, 1.953953e-08, -9.89246e-10, 4.371071e-08, 
    3.741167e-08, -1.045767e-07, -2.348935e-08, -7.69063e-09, 3.440559e-08, 
    -2.291637e-08, -1.806872e-08, 5.723248e-08, 1.599033e-08, 1.593611e-08, 
    4.67918e-09, -1.464715e-07, 5.859363e-08, -8.077683e-08, 1.219541e-07, 
    1.158738e-07, -1.359252e-07, 2.605526e-08, -6.75775e-08, -4.048445e-08, 
    1.951634e-08, -8.880846e-08, -1.781515e-08, -1.298205e-08, -1.797099e-08, 
    1.057117e-07, -1.666832e-07, 7.642427e-09, -6.507292e-08, -6.070665e-08, 
    3.934025e-08, -6.526903e-09, 3.671417e-09, -8.250893e-10, 5.75904e-08, 
    -3.86305e-08, -1.293921e-08, 5.5567e-08, -6.84355e-09, -2.551531e-09, 
    -6.291367e-08, -1.211794e-08, 2.913623e-09, -1.69868e-08, -5.399727e-09, 
    2.217644e-09, 1.399188e-08, -1.240732e-09, -1.195488e-09, -1.293849e-07,
  -1.448132e-08, 5.241361e-08, -2.879119e-09, -3.487571e-09, -2.669151e-08, 
    1.299179e-08, 6.744415e-08, 3.313687e-08, 3.315961e-08, -2.221782e-09, 
    -6.997436e-08, -1.093974e-08, 5.338359e-08, 1.455533e-09, -5.961112e-08, 
    -2.186562e-08, 3.346077e-09, 6.154153e-08, -6.044297e-08, -5.804884e-08, 
    8.260679e-08, 6.216521e-08, -4.652532e-08, -3.466687e-08, 6.867822e-10, 
    -4.461651e-08, 1.971068e-08, 3.842047e-09, -3.075832e-08, 1.274392e-07, 
    8.22032e-08, 1.152318e-08, 1.933915e-08, -1.583836e-07, -1.404393e-07, 
    -2.731497e-08, -3.008608e-08, 3.08807e-08, 1.038289e-07, 1.935252e-07, 
    -8.86994e-08, 3.39486e-08, -1.551325e-07, 6.931432e-08, -3.514458e-08, 
    -3.971979e-08, 1.09826e-08, 2.372656e-07, -3.854291e-08, -3.325667e-09, 
    5.976858e-09, -1.101008e-07, -8.077631e-09, -6.430833e-09, 1.012622e-08, 
    -2.889692e-09, 8.56777e-08, 1.898386e-07, 1.301078e-07, 1.010724e-08, 
    -6.478899e-09, -8.457653e-08, 5.419463e-08, -1.169412e-07, 2.055997e-08, 
    -4.286755e-08, 3.944058e-08, 1.677984e-08, -7.920221e-09, 3.819639e-08, 
    2.720105e-08, -4.697802e-08, -3.610705e-08, -1.950309e-08, 2.869826e-08, 
    -2.16445e-08, 1.650642e-08, 5.288456e-08, -9.039724e-09, 2.53259e-08, 
    -3.567266e-09, -9.672465e-08, 3.440027e-08, -6.956122e-08, -8.209213e-09, 
    -2.028276e-08, -1.477212e-07, -3.939249e-10, -9.943577e-08, -5.11501e-08, 
    -4.240121e-08, -7.372284e-08, -3.993227e-08, -7.457525e-08, 1.547289e-08, 
    1.573752e-07, -6.425815e-08, 7.020378e-08, -7.679648e-08, -7.076717e-08, 
    7.518679e-09, -2.570728e-08, 5.354153e-09, -2.627928e-09, 7.728306e-08, 
    -6.261405e-08, -3.142702e-08, 2.372951e-08, -2.411059e-08, -1.286787e-08, 
    -3.746015e-08, -7.909523e-08, 1.171543e-09, -3.212449e-09, 5.783556e-08, 
    3.543801e-09, 1.139662e-08, -2.255973e-09, -1.14423e-09, -4.314791e-08,
  -2.039332e-08, 7.948125e-08, -1.268012e-08, -5.538294e-08, -4.624411e-08, 
    -1.49027e-08, 3.454721e-08, 1.479123e-09, 2.919347e-08, -1.545453e-08, 
    -3.666213e-08, -3.277268e-08, 3.43137e-08, 2.961571e-08, -9.252852e-08, 
    3.132562e-08, 4.358719e-09, 2.101893e-08, -9.277397e-08, -2.565133e-08, 
    1.843665e-08, 9.013849e-08, -7.435887e-08, 7.615256e-09, 1.427689e-07, 
    2.04455e-08, 2.133612e-08, -1.98965e-08, -4.46143e-08, 1.378913e-07, 
    8.299418e-08, 2.079452e-08, 1.074756e-08, -1.367429e-07, -1.117716e-07, 
    -2.768201e-08, -2.721926e-08, 3.174679e-08, 1.064832e-07, 2.302791e-07, 
    -8.014126e-08, 2.833514e-08, -4.690565e-08, 8.946293e-08, -3.452277e-08, 
    -2.850919e-08, 5.674468e-08, 2.329728e-07, -3.115796e-08, 5.735501e-10, 
    6.922591e-09, -8.723754e-08, -4.666484e-08, 3.842273e-10, -8.821718e-09, 
    -8.939764e-10, 3.699967e-08, 1.732997e-07, 1.738755e-07, -1.602422e-08, 
    -2.911992e-08, 9.329011e-08, 7.807768e-08, -9.520312e-08, -6.450034e-09, 
    -4.454631e-08, 4.234954e-08, -7.369351e-09, -1.682128e-08, 2.354255e-08, 
    1.460722e-08, -5.243209e-08, -6.266094e-08, -2.840801e-08, 9.599972e-09, 
    -4.186035e-08, 2.887188e-08, 4.165537e-08, -1.760832e-08, 8.699345e-08, 
    -5.071399e-09, -7.531563e-08, 2.207872e-08, -7.810098e-08, 5.724752e-08, 
    -9.402169e-08, -4.368184e-08, -8.865925e-09, -1.069575e-07, 
    -2.172527e-08, -1.852461e-07, -6.72558e-08, -2.764614e-08, -1.394002e-07, 
    -5.227838e-08, 1.798504e-07, -7.848427e-09, 6.224133e-08, -7.053922e-08, 
    -4.284911e-08, 2.653343e-08, -3.19057e-07, 8.012663e-09, -3.38224e-09, 
    3.505653e-08, -9.266358e-08, -3.362305e-08, -1.126472e-08, -3.707345e-08, 
    -1.840471e-08, -3.183612e-08, -7.774355e-08, -7.104512e-08, 
    -7.391407e-09, 3.127803e-08, 3.066987e-09, 9.717184e-09, -2.464908e-09, 
    -1.051077e-09, 2.727808e-08,
  -5.348945e-07, 6.753788e-08, -2.060932e-08, -6.218949e-08, -2.974281e-08, 
    -4.366547e-08, -9.347849e-08, -9.904164e-08, 1.911548e-08, 1.412188e-07, 
    2.110073e-07, -2.185942e-08, 1.616678e-08, 3.022049e-07, -1.073875e-07, 
    6.195676e-08, 7.493441e-10, 7.652375e-09, -4.793323e-08, -3.448707e-08, 
    -1.992856e-08, 9.024092e-08, -5.60089e-08, 7.195484e-08, 2.27331e-08, 
    1.067852e-07, 2.958728e-08, -1.828511e-08, -2.928624e-08, 1.28256e-07, 
    4.83023e-08, 2.327801e-08, -1.409188e-08, -8.243211e-08, -4.63217e-10, 
    -4.289171e-08, -1.975687e-08, 3.208535e-08, 1.016275e-08, 2.27715e-07, 
    -6.599672e-08, 5.236228e-08, 2.09161e-09, 9.810663e-08, -5.549219e-08, 
    -3.267627e-08, 1.91657e-07, 1.849014e-07, -2.702406e-08, 3.249333e-09, 
    8.105218e-09, -8.929993e-08, -7.116671e-08, 4.443484e-09, -2.638291e-08, 
    -1.206502e-09, 2.700716e-08, 1.495411e-07, 7.327989e-08, -5.661774e-08, 
    2.427233e-07, 5.764883e-08, 9.104468e-08, -5.209749e-08, -1.951272e-08, 
    -4.072939e-08, 2.349651e-08, -9.511325e-09, -1.786867e-08, 4.025532e-08, 
    -8.33154e-10, -8.772889e-08, 6.128238e-08, -3.038366e-08, 7.833819e-09, 
    -2.752057e-08, 2.631465e-08, 2.465538e-08, -1.917668e-08, 7.412046e-08, 
    -2.550962e-09, -7.016418e-08, 3.316131e-09, -6.150555e-08, 1.218979e-08, 
    -1.494138e-07, 4.497394e-09, -8.599329e-09, -1.606212e-07, 3.089252e-08, 
    -8.658134e-08, -6.369829e-08, -6.798444e-09, -1.515898e-07, 
    -1.083914e-07, 1.163422e-07, -4.183804e-08, 6.960482e-08, -4.330246e-08, 
    -1.490822e-08, 1.481777e-08, 2.92109e-08, 7.216286e-09, -2.106532e-09, 
    -1.078905e-08, -1.03739e-07, -2.172368e-08, -3.625581e-08, -4.367399e-08, 
    -2.122175e-08, -2.817359e-08, -3.452948e-08, -9.769821e-08, 
    -6.355663e-10, 6.773064e-09, 1.251635e-09, 8.606719e-09, -2.541725e-09, 
    -8.847465e-10, -2.259259e-08,
  -1.519827e-06, -1.798679e-08, -3.210511e-08, -4.951204e-08, -6.219301e-08, 
    -1.436073e-07, -1.48072e-07, -1.19357e-07, -8.504287e-09, 8.233195e-08, 
    -9.887373e-08, 1.003485e-07, 4.442546e-08, 2.367716e-08, -4.247892e-08, 
    8.942207e-08, -1.055055e-08, 4.443689e-08, -2.916295e-08, -2.409087e-08, 
    -3.414135e-08, 5.37197e-08, -3.765859e-08, 1.646374e-07, 2.371013e-08, 
    2.348048e-07, 8.931863e-09, -1.263919e-08, -2.784628e-08, 1.034132e-07, 
    3.444194e-08, 1.159157e-08, -2.355392e-08, -4.542534e-08, 6.641875e-08, 
    -2.748078e-08, -2.446177e-09, 3.16323e-08, 4.849824e-09, 2.162361e-07, 
    -7.099938e-08, -1.174012e-07, 6.206491e-08, 9.985185e-08, -1.880079e-08, 
    -4.63869e-08, 1.787084e-07, 1.168904e-07, -8.856148e-09, 3.537032e-09, 
    9.214432e-09, -1.03296e-07, -8.330468e-08, 1.14588e-08, -3.996398e-08, 
    -1.077979e-09, 2.110136e-08, 1.0995e-08, -5.186433e-08, -7.743894e-08, 
    -7.316208e-08, -1.555321e-08, -1.278389e-07, -4.664614e-09, 
    -1.164688e-07, -3.608721e-08, 7.65624e-10, 7.388309e-08, -1.735185e-08, 
    6.477165e-08, -1.286679e-08, -8.773537e-08, 9.931853e-09, 5.794448e-09, 
    1.859583e-08, 1.834593e-08, 1.659406e-08, 3.974225e-08, -1.184407e-08, 
    -7.283518e-09, 3.243258e-09, -6.894825e-08, 1.993777e-08, -9.193496e-08, 
    -3.112444e-08, -1.22711e-07, -2.941903e-08, -7.573306e-09, -1.120297e-07, 
    7.346637e-08, -7.714056e-08, -7.01517e-08, -6.959823e-09, -1.206337e-07, 
    -1.521204e-08, -1.5258e-07, -5.26764e-08, -2.271264e-08, -2.563223e-08, 
    -6.922516e-09, 6.818829e-08, 2.378863e-07, -4.56062e-08, 5.375895e-10, 
    3.149881e-08, -1.056432e-07, -3.973759e-08, -6.864587e-08, -4.804468e-08, 
    -2.209566e-08, -2.62873e-08, -1.184543e-08, -2.476753e-08, 7.229914e-10, 
    3.597791e-09, -3.954142e-10, 7.655117e-09, -2.797002e-09, -8.540226e-10, 
    -7.272257e-08,
  -1.390905e-06, -1.005685e-07, -4.388062e-08, -1.145188e-07, -1.838885e-07, 
    -1.765596e-07, -8.54094e-08, -7.121139e-08, -4.676622e-09, -1.111214e-07, 
    -9.529447e-08, 1.438457e-08, 3.210159e-07, -8.700943e-08, 7.233734e-08, 
    1.138494e-07, -8.31252e-09, 1.358967e-08, 3.188457e-08, -3.506068e-08, 
    -1.131298e-08, 7.838707e-10, 1.643839e-07, 2.936304e-09, -1.28878e-07, 
    1.158493e-07, -1.367994e-08, -6.649884e-09, -1.447052e-08, 9.434575e-08, 
    4.92538e-08, -2.141815e-08, -1.350668e-08, -5.812774e-08, 6.049993e-08, 
    -2.294473e-08, 1.230428e-08, 3.154396e-08, -2.68642e-10, 1.88441e-07, 
    -9.472335e-08, 2.81243e-08, 7.467571e-08, 8.350518e-08, 4.684091e-08, 
    -7.159895e-08, 2.065385e-07, 4.519319e-08, -2.948855e-09, 2.790152e-09, 
    1.075084e-08, 5.594893e-08, -1.323233e-07, 2.652318e-08, -5.550637e-08, 
    -9.252403e-10, 1.354658e-08, -5.050003e-08, -1.438778e-09, -7.867588e-08, 
    -1.594559e-07, -3.354035e-08, -1.883677e-08, 2.219925e-08, -1.722983e-07, 
    -3.580431e-08, -1.083595e-08, 8.559209e-08, -2.12035e-08, 7.351946e-08, 
    2.946081e-09, -8.079621e-08, -6.307914e-09, 7.756e-08, 5.730378e-09, 
    3.418131e-08, -5.077482e-09, 1.528065e-08, 5.340414e-09, -9.206019e-08, 
    1.362162e-08, -6.528643e-08, -4.470678e-09, -9.484586e-08, -5.330844e-08, 
    -8.286634e-08, -6.26419e-08, -1.411388e-08, -4.815919e-08, 9.887833e-08, 
    -6.404025e-08, -7.208714e-08, -5.660894e-09, -6.921262e-08, 
    -2.274624e-08, -6.020081e-08, -4.918857e-08, 1.010869e-08, -2.214085e-08, 
    -4.930007e-08, 1.407575e-07, 1.414884e-07, -9.871997e-08, 3.199084e-09, 
    3.729133e-08, -8.763834e-08, -7.743165e-08, -9.824237e-08, -5.370941e-08, 
    -2.259003e-08, -2.47029e-08, -7.007998e-09, 3.301807e-09, 1.084572e-09, 
    2.029651e-09, -1.267142e-09, 6.059366e-09, -2.482672e-09, -8.587904e-10, 
    -1.027056e-07,
  -4.429431e-07, 1.096794e-08, -1.490321e-07, -3.240356e-07, -1.580277e-07, 
    -4.288802e-08, -4.611695e-08, -1.054698e-07, -2.01502e-08, -1.068631e-07, 
    8.876782e-09, 1.281262e-08, -2.206946e-08, -1.03178e-07, 9.104247e-08, 
    1.053453e-07, -3.397835e-08, 8.292432e-09, 7.073767e-08, 5.624111e-08, 
    -2.618924e-08, -7.425342e-09, 1.004995e-07, -1.747151e-08, -6.009668e-08, 
    -1.296507e-08, -1.647254e-08, 4.105232e-10, -2.179399e-08, 9.837356e-08, 
    4.632295e-08, -1.439003e-08, 9.307996e-09, -6.371329e-08, 8.931465e-09, 
    -1.339902e-08, -5.736499e-08, 3.133728e-08, -1.15233e-09, 1.475149e-07, 
    -1.085291e-07, 8.895643e-08, -1.801141e-09, 8.767354e-08, 6.187713e-08, 
    -8.150016e-08, 2.212862e-07, -3.88161e-09, -1.350602e-08, 2.469022e-09, 
    1.296648e-08, -1.097236e-07, -1.008137e-07, 3.605055e-08, -5.447128e-08, 
    1.065075e-09, 4.072012e-08, -9.167798e-08, -4.97743e-09, -6.633898e-08, 
    -9.021335e-08, -3.002697e-08, 4.19335e-08, 2.747709e-08, -1.900142e-07, 
    -4.024048e-08, -7.403401e-09, 6.977189e-08, -2.008517e-08, 6.510902e-08, 
    2.484762e-08, -4.746164e-08, -5.594814e-08, 1.167291e-08, 4.540347e-09, 
    1.786702e-08, 1.927543e-08, 1.483937e-08, 1.229797e-08, -7.081178e-08, 
    3.654827e-08, -2.712963e-08, 4.615288e-09, -5.992104e-08, -5.92762e-08, 
    -1.138072e-07, 6.974119e-09, -4.241849e-08, 3.402739e-09, 1.202146e-07, 
    -7.448875e-08, -6.640958e-08, 7.74719e-10, -3.119089e-08, -2.688455e-08, 
    -3.554469e-08, 6.274465e-08, 8.276072e-08, -2.72496e-08, -3.456869e-08, 
    1.067486e-07, 6.331416e-08, -3.637839e-08, 5.474114e-09, 1.515559e-09, 
    -6.379207e-08, -1.070249e-07, -1.160374e-07, -5.170045e-08, 
    -1.703518e-08, -2.533579e-08, -4.45732e-09, 6.830192e-09, 1.320927e-09, 
    5.461516e-10, -1.652916e-09, 6.006118e-09, -2.199894e-09, -7.12852e-10, 
    7.046742e-08,
  -1.767506e-08, 7.916929e-07, -1.339067e-07, -2.411697e-07, -1.576945e-07, 
    1.707036e-08, -1.6304e-08, -3.678286e-08, 4.931809e-08, -1.978441e-08, 
    1.033897e-08, 8.599551e-08, 2.132932e-07, -2.018936e-08, 1.328345e-08, 
    1.167823e-07, -4.771838e-08, 2.828159e-08, 5.906145e-08, 5.409544e-08, 
    -5.649667e-10, -8.057839e-09, 4.470081e-08, -2.491873e-08, -2.279484e-08, 
    -2.886003e-08, 1.306768e-08, 6.643461e-09, 4.080567e-08, 2.053173e-07, 
    5.747785e-08, -3.438953e-08, 5.181903e-09, 2.544567e-08, -7.547845e-08, 
    -7.677443e-09, -6.196084e-08, 3.001452e-08, 1.553946e-08, 1.113285e-07, 
    -1.010724e-07, 6.980105e-08, -1.206604e-08, 7.208739e-08, 7.310547e-08, 
    -8.518754e-08, 2.106089e-07, -1.25404e-08, -1.9786e-08, 1.878362e-09, 
    1.479316e-08, -1.276268e-07, -4.506695e-08, 3.974006e-08, -4.932316e-08, 
    2.159311e-09, -5.518535e-08, -9.995501e-08, -7.163713e-09, -7.58186e-08, 
    -4.038833e-08, 1.881773e-08, -1.902123e-07, 2.914027e-08, -1.67737e-07, 
    -2.142764e-08, 5.936101e-09, 4.688746e-08, -2.025985e-08, 5.239104e-08, 
    -4.659836e-08, -1.21874e-08, -2.524227e-07, -1.326765e-08, 4.785928e-09, 
    4.364495e-09, 8.102268e-08, 3.841251e-08, 1.566794e-08, -1.32914e-07, 
    3.958991e-08, 4.355923e-09, 1.392897e-08, 6.766396e-08, -1.282154e-08, 
    -1.846658e-07, 1.127615e-07, -1.057853e-07, 5.186804e-08, 1.391275e-07, 
    2.184612e-08, -3.822005e-08, -7.705694e-10, -1.104432e-08, 6.501182e-10, 
    -2.362218e-08, 3.460892e-08, 6.919169e-08, -2.989367e-08, -1.055326e-08, 
    4.192435e-08, -4.042931e-09, -1.439473e-08, 6.814787e-09, 5.911176e-08, 
    -6.103272e-08, -1.282817e-07, -1.262528e-07, -4.288671e-08, 
    -1.386906e-08, -2.650717e-08, -3.543335e-09, 8.326253e-09, 1.725596e-09, 
    -1.025171e-09, -1.638239e-09, 9.599006e-09, -2.238615e-09, -7.575238e-10, 
    4.320157e-09,
  1.988499e-07, 2.187954e-07, 2.359377e-08, -8.494112e-09, -6.832715e-08, 
    3.260959e-08, -1.09743e-08, -2.856518e-08, 2.92797e-08, -1.356977e-08, 
    6.510845e-08, 8.385427e-09, -9.052656e-09, 8.063807e-10, -8.557436e-09, 
    1.568275e-07, -7.769422e-08, 2.098847e-08, 3.447735e-08, -6.498135e-08, 
    -1.282922e-08, -3.461423e-09, 1.681747e-08, -2.93802e-08, 1.154376e-09, 
    -3.355717e-08, -1.135788e-08, 1.38449e-08, 5.707852e-08, 3.146619e-07, 
    9.394807e-08, 8.4833e-08, -3.418518e-08, -5.947004e-08, -1.170213e-08, 
    4.442938e-08, -5.315724e-08, 2.688164e-08, 7.909648e-08, 8.760802e-08, 
    -6.682023e-08, 2.473973e-08, -1.479785e-08, 3.918183e-08, 7.272922e-08, 
    -8.398547e-08, 1.695885e-07, -1.288424e-08, -1.941432e-08, 1.18925e-09, 
    1.641862e-08, -1.154789e-07, -7.322984e-08, 3.578512e-08, -4.61023e-08, 
    3.154412e-09, -1.252639e-07, -1.054198e-07, -8.991272e-09, -8.161049e-08, 
    -3.967534e-08, 2.629554e-08, 1.095954e-07, 4.636522e-08, -7.288259e-09, 
    -3.857849e-09, 1.815783e-08, 2.535955e-08, -3.063519e-08, 3.149137e-08, 
    -3.569551e-08, -9.562541e-09, -3.225625e-08, -2.387424e-11, 4.849745e-09, 
    -1.13813e-08, 5.401702e-09, 2.795053e-08, 3.615571e-08, -3.167165e-07, 
    5.975596e-08, 1.585502e-08, 1.056003e-08, -6.06758e-09, 1.563785e-08, 
    -2.414e-07, -4.84373e-08, -1.311879e-07, 7.545113e-08, 1.535475e-07, 
    3.464731e-08, -1.044264e-08, -5.106813e-10, 1.367083e-08, -1.679723e-08, 
    -1.851856e-08, 5.230495e-08, 1.167002e-07, -3.0249e-08, 6.481923e-09, 
    -4.325989e-08, -2.708938e-08, 3.542831e-08, 7.8659e-09, 6.310984e-08, 
    -5.557649e-08, -1.398065e-07, -1.32971e-07, -3.563684e-08, -1.157468e-08, 
    -2.79307e-08, -2.946422e-09, 9.624273e-09, 2.270212e-09, -3.469722e-09, 
    -3.820673e-10, 1.351012e-09, -3.717361e-09, -9.56959e-10, 3.759965e-09,
  2.397188e-07, 1.784249e-07, 1.518526e-08, 5.727998e-09, 3.770128e-08, 
    -5.431275e-09, 1.213266e-09, 5.763957e-08, 1.577325e-08, 2.006414e-08, 
    9.356427e-10, 4.20107e-09, 5.029278e-09, 1.844637e-08, -8.262759e-09, 
    2.095624e-07, -6.661632e-08, -4.918832e-09, 2.880024e-08, -7.289236e-08, 
    -1.411479e-08, -2.094339e-09, 1.017497e-09, -3.075968e-08, 1.233991e-08, 
    -3.511104e-08, -3.757577e-08, 1.82331e-09, 3.856462e-08, 3.00691e-07, 
    1.962394e-08, 6.632979e-08, 4.152253e-08, -1.751396e-07, -1.258343e-08, 
    1.027993e-07, -4.47266e-08, 2.237866e-08, 4.510423e-08, 7.214575e-08, 
    -2.57989e-08, 1.61848e-08, -1.638222e-08, 2.359474e-08, 4.934509e-08, 
    -9.10876e-08, 1.202496e-07, -1.637457e-08, -2.228344e-08, -2.130207e-11, 
    1.764204e-08, -1.253907e-07, -6.336727e-08, 3.558373e-08, -4.182262e-08, 
    1.737874e-09, -1.529776e-07, -1.082525e-07, -1.030813e-08, -1.87907e-08, 
    -2.787431e-08, 2.757645e-08, 9.151427e-08, 6.841381e-08, -5.699392e-08, 
    3.398907e-08, -4.058586e-08, 3.527066e-08, -1.441015e-08, 1.044884e-08, 
    4.218919e-10, 1.31962e-08, 5.1906e-09, -7.410108e-09, 4.683592e-09, 
    -1.881949e-08, -4.978062e-10, 2.437525e-08, 4.680622e-08, -9.669884e-08, 
    5.716174e-08, 2.053986e-08, 7.930225e-09, -1.220815e-08, 2.110335e-08, 
    -1.503669e-07, -6.68158e-08, -1.889657e-08, 1.042696e-07, 1.575849e-07, 
    3.404955e-08, -1.314015e-08, -1.363674e-10, 4.517736e-08, -2.332802e-07, 
    -1.756951e-08, 5.029433e-08, 2.257874e-07, -2.894751e-08, 3.196944e-08, 
    -1.322162e-07, -3.949192e-08, 3.589532e-08, 8.801635e-09, 7.109463e-08, 
    -3.847902e-08, -1.700008e-07, -1.379889e-07, -3.197135e-08, 
    -1.139745e-08, -2.925253e-08, -2.764523e-09, 1.061449e-08, 2.872525e-09, 
    -6.575306e-09, 1.112005e-09, 3.689067e-09, -1.855586e-09, -1.012879e-09, 
    5.014954e-09,
  2.491704e-07, 1.664694e-07, 1.033357e-08, 5.775632e-09, 4.550554e-08, 
    1.8984e-08, 2.927266e-08, 5.559082e-08, 2.207469e-08, 2.808838e-08, 
    3.34262e-09, 4.779622e-09, 9.396786e-09, 2.154786e-08, -8.129632e-09, 
    2.248949e-07, -4.781159e-08, 7.961546e-09, -3.155462e-08, -7.590779e-08, 
    -1.464934e-08, -1.174726e-09, -5.851462e-09, -3.118862e-08, 1.807916e-08, 
    -3.591697e-08, -3.782566e-08, -5.948755e-08, -1.068306e-07, 1.949638e-08, 
    2.355557e-08, 9.786686e-08, 4.547974e-08, -1.77935e-07, -1.279523e-08, 
    1.047956e-07, -3.804094e-08, 1.788733e-08, 1.929868e-08, 6.239154e-08, 
    -4.106066e-08, 1.175408e-08, -1.689006e-08, 2.338638e-08, 1.389365e-07, 
    -8.301606e-08, 5.833272e-08, -2.267979e-08, -1.793294e-08, -6.735377e-10, 
    1.864342e-08, -1.240765e-07, -5.645446e-08, 3.765906e-08, -3.240381e-08, 
    2.425963e-09, -1.846287e-07, -1.096254e-07, -1.131512e-08, 1.126034e-07, 
    -1.973365e-08, 2.810827e-08, 9.78705e-08, 7.908291e-08, -7.359713e-08, 
    1.573864e-07, -7.152232e-08, 7.758149e-08, -1.36647e-08, 9.525934e-09, 
    -2.431875e-09, -1.298019e-08, 1.679132e-08, -8.534585e-09, 4.48923e-09, 
    -3.442563e-08, -2.38191e-09, 2.124855e-08, 4.923042e-08, -3.647381e-08, 
    1.402572e-08, 1.434107e-08, 6.184678e-09, -1.368028e-08, 9.572204e-09, 
    -7.181063e-08, -6.427581e-08, 3.356854e-08, 1.06604e-07, 1.593754e-07, 
    3.376874e-08, -2.018937e-08, 2.552554e-10, 6.68453e-08, -8.707468e-08, 
    -1.630571e-08, 5.462182e-08, -6.011339e-08, -1.867681e-08, 2.8571e-08, 
    -9.801715e-08, -4.681934e-08, 3.222703e-08, 9.212179e-09, 7.08269e-11, 
    -2.822367e-08, -1.891262e-07, -1.349573e-07, -3.238165e-08, 
    -1.229159e-08, -2.974753e-08, -2.429147e-09, 1.159356e-08, 3.425384e-09, 
    -6.61521e-09, 6.14009e-09, 9.636665e-10, -1.536584e-09, -8.881855e-10, 
    5.482661e-09,
  2.480789e-07, 1.601906e-07, 8.784696e-09, 3.901505e-09, 4.941796e-08, 
    3.149728e-08, 3.300534e-08, 5.536572e-08, 2.329773e-08, 3.279138e-08, 
    4.278036e-10, 4.41662e-09, 1.078831e-08, 2.006038e-08, -8.006054e-09, 
    2.184156e-07, -9.204245e-09, 1.682685e-08, -4.754749e-08, -7.731444e-08, 
    -1.484318e-08, 1.115609e-09, -5.303718e-09, -3.160119e-08, 2.101785e-08, 
    -3.567925e-08, -2.653883e-08, -4.943331e-09, -1.099198e-07, 
    -3.361674e-08, 2.411753e-08, 1.298199e-07, -1.262994e-07, 1.45238e-07, 
    -1.284843e-08, 2.746276e-08, -3.161226e-08, 1.319123e-08, 5.744459e-08, 
    5.80094e-08, 5.326662e-09, 9.405881e-09, -1.875719e-08, 1.524457e-08, 
    9.026587e-08, -8.351356e-08, 2.221481e-08, -2.922624e-08, -1.667052e-08, 
    -1.063619e-09, 1.936493e-08, -1.226912e-07, -5.327924e-08, 3.826697e-08, 
    -1.704067e-08, 5.848051e-10, -1.881664e-07, -1.113755e-07, -1.226598e-08, 
    2.3765e-08, -1.786611e-08, 2.82688e-08, 9.973996e-08, 8.830243e-08, 
    -3.255054e-08, 1.894955e-08, -2.225465e-08, -6.177061e-09, 1.470585e-08, 
    -3.293246e-08, 4.083631e-10, -3.597438e-08, 2.088564e-08, -8.953634e-09, 
    3.992319e-09, -3.247908e-08, -3.702837e-09, 1.721421e-08, 4.177884e-08, 
    -1.154217e-08, -2.347696e-08, 7.935959e-09, 5.612094e-09, -1.411217e-08, 
    6.671144e-09, -1.592125e-07, -6.809626e-08, 2.609465e-08, 1.000194e-07, 
    1.585232e-07, 3.353296e-08, -3.103712e-08, 9.416112e-10, 7.405865e-08, 
    8.487973e-09, -1.559255e-08, 5.888607e-08, -7.389031e-08, -1.326623e-08, 
    2.552181e-08, -1.263724e-07, -4.938041e-08, 2.74372e-08, 8.987669e-09, 
    2.677757e-08, 1.292847e-08, -1.882994e-07, -1.289189e-07, -3.42061e-08, 
    -1.309013e-08, -2.871332e-08, -2.365482e-09, 1.20333e-08, 4.333288e-09, 
    1.14585e-09, 1.21305e-09, 4.515101e-09, -1.173944e-09, -7.033805e-10, 
    5.79621e-09,
  2.477252e-07, 1.558712e-07, 8.275492e-09, 3.492005e-09, 5.128516e-08, 
    3.176365e-08, 3.530204e-08, 5.469474e-08, 2.339732e-08, 3.485354e-08, 
    -4.303956e-09, 5.528591e-09, 1.125045e-08, 2.102217e-08, -7.885205e-09, 
    1.975896e-07, 1.33206e-08, 1.832825e-08, -5.766233e-08, -7.805022e-08, 
    -1.507397e-08, -2.310344e-09, -1.219519e-09, -3.269793e-08, 2.316642e-08, 
    -3.538582e-08, -3.619573e-08, 5.310312e-09, -1.127084e-07, -6.179516e-08, 
    4.098808e-08, 5.863558e-08, -1.041921e-07, 2.543595e-08, -1.286378e-08, 
    2.22883e-09, -2.559428e-08, 7.114991e-09, -7.63373e-09, 5.755282e-08, 
    4.280073e-08, 7.950575e-09, -1.902009e-08, 1.669415e-08, 3.733624e-08, 
    -8.432437e-08, -1.518231e-09, -3.373214e-08, -1.614606e-08, 
    -1.670294e-09, 1.967641e-08, -1.211719e-07, -5.279272e-08, 4.064736e-08, 
    -9.175514e-09, 2.441993e-10, -1.62893e-07, -1.122723e-07, -1.341918e-08, 
    -1.728033e-08, -1.734679e-08, 2.836703e-08, 1.029447e-07, 1.044729e-07, 
    -1.93472e-08, -1.099784e-08, -3.064906e-08, -6.045764e-08, -1.366175e-08, 
    -3.621597e-08, 2.424315e-08, -3.677553e-08, 2.257377e-08, -9.189534e-09, 
    3.366324e-09, -1.528224e-08, -3.872671e-09, 1.759588e-08, 1.708287e-08, 
    -8.728762e-09, -4.830918e-08, 4.433893e-09, 2.86002e-09, -1.423143e-08, 
    5.770744e-09, -9.767723e-08, -7.128301e-08, 2.475338e-08, 9.114046e-08, 
    1.564777e-07, 3.292632e-08, -4.194769e-08, 1.752738e-09, 6.787955e-08, 
    3.601201e-08, -1.5347e-08, 6.204407e-08, -8.118104e-08, -9.506152e-09, 
    2.405452e-08, -1.121218e-07, -4.895207e-08, 2.864763e-08, 9.717617e-09, 
    2.634476e-08, 1.468993e-08, -1.672109e-07, -1.279199e-07, -3.670118e-08, 
    -1.370745e-08, -2.560625e-08, -2.059323e-09, 1.192234e-08, 4.910135e-09, 
    2.388413e-08, 2.077511e-10, 4.078245e-09, -1.648662e-09, -6.635403e-10, 
    6.102255e-09,
  2.471668e-07, 1.517999e-07, 8.75491e-09, 2.664933e-09, 5.246932e-08, 
    3.361947e-08, 3.636649e-08, 5.370759e-08, 2.294632e-08, 3.557659e-08, 
    -4.965386e-09, 5.570314e-09, 1.144292e-08, 2.200034e-08, -7.946142e-09, 
    1.955688e-07, 2.199747e-08, 2.052934e-08, -6.640279e-08, -7.83956e-08, 
    -1.531976e-08, -4.57112e-09, 1.765329e-09, -3.296873e-08, 2.459092e-08, 
    -3.495518e-08, -3.803757e-08, 2.689035e-08, -1.15788e-07, -7.685651e-08, 
    5.426182e-08, 6.260063e-08, -4.285675e-08, 4.54537e-08, -1.316539e-08, 
    2.493664e-08, -2.019137e-08, 2.496321e-09, 2.324509e-08, 5.937897e-08, 
    5.503605e-08, 6.719802e-09, -1.953828e-08, 1.283284e-08, 1.744286e-08, 
    -8.548477e-08, -2.584738e-08, -3.764617e-08, -1.597596e-08, 
    -1.950418e-09, 1.965391e-08, -1.20043e-07, -5.383515e-08, 4.206204e-08, 
    -1.154227e-08, 1.191779e-09, -1.816101e-07, -1.121553e-07, -1.490735e-08, 
    -3.522484e-08, -1.660169e-08, 2.768888e-08, 1.043106e-07, 1.17602e-07, 
    -1.374681e-08, -1.78602e-08, -6.262894e-09, -6.925745e-08, -9.86654e-09, 
    -4.201684e-08, 2.333275e-08, -5.473612e-08, 2.335628e-08, -9.301743e-09, 
    2.564569e-09, -1.374292e-08, -3.675552e-09, 1.783738e-08, 4.677585e-09, 
    -4.173899e-09, -2.678661e-08, 9.564047e-10, 6.189737e-09, -1.385638e-08, 
    4.872049e-09, -7.410631e-08, -7.309734e-08, 2.486786e-08, 8.402719e-08, 
    1.544877e-07, 3.246305e-08, -4.47528e-08, 2.350845e-09, 5.521342e-08, 
    4.432775e-08, -1.486116e-08, 6.447844e-08, -8.151039e-08, -7.262202e-09, 
    2.47481e-08, -1.003976e-07, -4.801023e-08, 2.570074e-08, 9.311933e-09, 
    2.607158e-08, 1.623596e-08, -1.356561e-07, -1.356602e-07, -4.175172e-08, 
    -1.33939e-08, -2.099659e-08, -7.613608e-10, 1.141666e-08, 4.768253e-09, 
    5.522975e-08, -1.143667e-09, 9.921251e-09, -9.946817e-10, -7.257981e-10, 
    5.782908e-09,
  2.459574e-07, 1.471799e-07, 8.013217e-09, 2.051138e-09, 5.375489e-08, 
    3.485184e-08, 3.708237e-08, 5.224501e-08, 2.202728e-08, 3.785544e-08, 
    -5.568722e-09, 5.077709e-09, 1.251885e-08, 2.236914e-08, -8.119969e-09, 
    1.921916e-07, 2.484213e-08, 2.150989e-08, -7.280494e-08, -7.891913e-08, 
    -1.546266e-08, -5.725724e-09, 1.746912e-09, -3.298112e-08, 2.495585e-08, 
    -3.434809e-08, -3.93668e-08, 3.635807e-08, -1.184983e-07, -8.434699e-08, 
    6.060054e-08, 5.641368e-08, -3.557193e-08, 1.035708e-07, -1.372712e-08, 
    2.952936e-08, -1.601404e-08, 2.305484e-09, 5.041795e-08, 5.924095e-08, 
    3.749938e-08, 5.6217e-09, -2.058295e-08, 1.103034e-08, 7.267431e-09, 
    -8.599875e-08, -4.645017e-08, -4.053746e-08, -1.631306e-08, 
    -2.131763e-09, 1.966819e-08, -1.188382e-07, -5.551858e-08, 4.994681e-08, 
    -2.625788e-08, -3.067271e-10, -1.951856e-07, -1.110482e-07, 
    -1.695831e-08, -4.211002e-08, -1.550632e-08, 2.636114e-08, 1.037191e-07, 
    1.248404e-07, -1.179874e-08, -2.041691e-08, -3.037337e-08, -8.328084e-08, 
    -1.643912e-08, -4.367701e-08, 1.653996e-08, -3.951232e-08, 2.305057e-08, 
    -9.140649e-09, 1.455806e-09, 1.359513e-08, -3.790461e-09, 2.02142e-08, 
    -2.536297e-09, -2.342858e-09, -1.926816e-08, -2.313435e-09, 1.422831e-08, 
    -1.287754e-08, 7.482868e-09, -6.991922e-08, -7.320102e-08, 2.477327e-08, 
    8.210311e-08, 1.521611e-07, 3.128412e-08, -4.53753e-08, 2.602235e-09, 
    4.308261e-08, 4.777883e-08, -1.4851e-08, 6.513812e-08, -8.536176e-08, 
    -6.511755e-09, 2.639936e-08, -9.606106e-08, -4.716745e-08, 2.315544e-08, 
    8.886715e-09, 2.632476e-08, 1.759361e-08, -8.12347e-08, -1.471064e-07, 
    -4.751723e-08, -1.219814e-08, -1.662909e-08, 2.315574e-09, 1.071203e-08, 
    5.052016e-09, 5.144511e-08, 7.230255e-10, 1.683496e-08, -1.290609e-09, 
    -2.153975e-09, 5.606125e-09,
  2.446715e-07, 1.409354e-07, 7.981043e-09, 4.039634e-09, 5.52235e-08, 
    3.636842e-08, 3.74198e-08, 4.997401e-08, 2.037314e-08, 3.775222e-08, 
    -5.803486e-09, 3.354216e-09, 1.315721e-08, 2.226659e-08, -8.431471e-09, 
    1.878223e-07, 2.418506e-08, 2.201523e-08, -7.92306e-08, -7.949313e-08, 
    -1.567264e-08, -6.072582e-09, 1.357307e-09, -3.276284e-08, 2.51116e-08, 
    -3.331138e-08, -3.887078e-08, 4.226126e-08, -1.205593e-07, -8.758275e-08, 
    6.037124e-08, 5.092932e-08, -3.33855e-08, 3.683282e-07, -1.546255e-08, 
    3.623654e-08, -1.402653e-08, 1.787541e-09, 7.484005e-08, 5.928327e-08, 
    1.887679e-08, 4.739945e-09, -2.221046e-08, 4.382487e-09, -1.958824e-10, 
    -8.866209e-08, -6.656467e-08, -4.227678e-08, -1.565704e-08, 
    -4.437616e-09, 2.019004e-08, -1.173019e-07, -5.73632e-08, 4.630829e-08, 
    -4.815057e-08, -5.856123e-09, -2.067601e-07, -1.09527e-07, -2.009093e-08, 
    -4.466618e-08, -1.403271e-08, 2.408171e-08, 1.003068e-07, 1.305789e-07, 
    -1.331271e-08, -2.222919e-08, -3.755486e-08, -9.547e-08, -2.842251e-08, 
    -4.412573e-08, 1.065291e-08, -4.142771e-08, 2.185652e-08, -9.176347e-09, 
    -2.78007e-10, 8.832785e-09, -3.260112e-09, 2.131901e-08, -3.367493e-09, 
    -1.911644e-09, -1.549699e-08, -5.080331e-09, 2.364163e-08, -1.166893e-08, 
    9.615178e-09, -7.440542e-08, -7.451638e-08, 2.435229e-08, 7.696579e-08, 
    1.483216e-07, 3.089974e-08, -4.289516e-08, 2.667633e-09, 3.390284e-08, 
    4.409935e-08, -1.548618e-08, 6.739567e-08, -8.575989e-08, -6.096116e-09, 
    2.728696e-08, -1.009469e-07, -4.612041e-08, 2.695682e-08, 8.489735e-09, 
    2.804461e-08, 1.924695e-08, 5.015715e-08, -1.556363e-07, -5.19176e-08, 
    -1.478566e-08, -1.643821e-08, 3.457103e-09, 1.012654e-08, 4.617164e-09, 
    3.208754e-08, 2.944944e-10, 3.251247e-08, 3.33079e-09, -4.496719e-09, 
    5.777224e-09,
  2.431686e-07, 1.282836e-07, 9.922076e-09, 5.202935e-09, 5.744988e-08, 
    3.922258e-08, 3.737722e-08, 4.493319e-08, 1.634004e-08, 3.573899e-08, 
    -5.903928e-09, 2.590525e-09, 1.301902e-08, 2.126291e-08, -9.122857e-09, 
    1.796783e-07, 2.212322e-08, 2.206849e-08, -7.991183e-08, -7.977684e-08, 
    -1.616996e-08, -6.89721e-09, 4.902745e-10, -3.197141e-08, 2.554901e-08, 
    -3.095948e-08, -4.130385e-08, 4.66801e-08, -1.224113e-07, -8.817773e-08, 
    5.678447e-08, 4.912937e-08, -3.241843e-08, 5.625297e-07, -1.931897e-08, 
    4.802047e-08, -1.754751e-08, 1.647223e-09, 3.78306e-08, 5.936742e-08, 
    4.349555e-09, 4.216247e-09, -2.562862e-08, 3.562548e-09, -4.264109e-09, 
    -9.102172e-08, -8.980743e-08, -4.3451e-08, -1.458146e-08, -8.591698e-09, 
    2.048937e-08, -1.14269e-07, -5.93299e-08, 4.522375e-08, -9.03739e-08, 
    -1.131292e-08, -1.865009e-07, -1.011697e-07, -2.606595e-08, 
    -4.698391e-08, -1.114353e-08, 2.030794e-08, 9.177558e-08, 1.320317e-07, 
    -1.5439e-08, -2.469238e-08, -3.940539e-08, -9.873912e-08, -3.289875e-08, 
    -4.363284e-08, 8.125028e-09, 1.405539e-08, 1.924928e-08, -9.271446e-09, 
    -4.015568e-09, -1.460165e-08, -1.457764e-09, 1.951994e-08, 7.626275e-09, 
    -2.223089e-09, -1.275839e-08, -7.256425e-09, 3.332366e-08, -9.153666e-09, 
    1.059294e-08, -6.729971e-08, -6.627789e-08, 2.318285e-08, 5.945279e-08, 
    1.474314e-07, 3.042459e-08, -3.857546e-08, 2.144503e-09, 2.615494e-08, 
    4.215866e-08, -1.758788e-08, 6.170732e-08, -8.384899e-08, -6.405514e-09, 
    2.731527e-08, -9.568697e-08, -4.498405e-08, 2.562794e-08, 8.021573e-09, 
    2.791563e-08, 2.280166e-08, 9.185857e-08, -1.607561e-07, -5.465421e-08, 
    -1.830932e-08, -1.840516e-08, 1.736623e-09, 1.217046e-08, 5.506479e-09, 
    2.776557e-08, 3.916625e-10, 6.93187e-08, 2.748209e-09, 8.678484e-09, 
    5.96259e-09,
  1.866098e-13, 4.056981e-13, 5.056766e-13, 5.601754e-13, 4.039193e-13, 
    1.272984e-13, -1.685365e-13, -2.14592e-13, 1.011997e-12, 3.684174e-13, 
    1.268585e-13, -3.98565e-13, 5.809993e-14, 1.756013e-14, -9.669973e-14, 
    -3.450422e-13, -1.686862e-12, -2.651818e-13, -2.01976e-13, -1.094683e-12, 
    -4.27087e-12, -8.743089e-13, 8.559743e-13, -7.555373e-13, -2.503275e-13, 
    1.05067e-13, 1.869724e-13, -3.978916e-14, 5.277076e-14, -1.229925e-13, 
    1.965481e-14, -1.346808e-13, 1.603248e-13, 2.755549e-14, 6.008798e-13, 
    -9.630363e-14, 3.538837e-14, 3.980314e-12, 3.511096e-13, 1.434161e-13, 
    1.706126e-12, -3.584497e-13, 7.659602e-14, -1.185933e-12, 2.030331e-13, 
    6.397828e-13, 1.052742e-12, 6.670329e-13, -1.867945e-12, 6.764283e-13, 
    5.219363e-13, 3.599429e-14, 4.126184e-13, -6.044502e-13, -1.131494e-13, 
    -1.631052e-12, -2.253458e-13, -4.566703e-13, 1.590062e-13, 1.545807e-12, 
    1.020666e-12, -3.915039e-13, 2.535699e-13, -5.9673e-13, -2.62125e-13, 
    -3.34667e-13, 7.433749e-13, -7.015332e-14, -8.082646e-14, 1.438239e-13, 
    7.700618e-14, 1.142257e-14, 8.807946e-14, 2.901897e-13, 6.692874e-13, 
    -5.333196e-14, 5.337515e-13, -1.230985e-12, -9.003271e-13, -2.567582e-13, 
    -3.287933e-13, 4.340541e-13, 1.690598e-13, -2.028826e-13, 7.596207e-13, 
    1.828115e-13, -3.429508e-13, -3.698852e-13, 7.243173e-14, 5.711753e-13, 
    1.151821e-13, 8.574951e-13, 5.024078e-13, 7.674461e-13, -3.819263e-14, 
    -3.939094e-13, -1.994388e-13, -4.440342e-13, -1.413801e-13, 
    -7.397398e-13, -6.746465e-13, 4.214286e-13, -5.145562e-13, 1.359503e-12, 
    5.92554e-14, 8.591417e-14, 4.08926e-13, -2.722936e-13, -7.666975e-13, 
    -5.232928e-13, -2.970424e-13, -8.823846e-14, -4.890319e-14, 
    -7.036743e-15, 5.334254e-13, -8.956529e-12, 1.116097e-12, -3.703339e-13, 
    -1.369756e-12, -1.157827e-13,
  -1.00131e-13, -1.230275e-13, -8.021354e-14, -4.234256e-14, -1.418647e-15, 
    4.698282e-14, 7.039488e-14, 9.391984e-14, 2.439967e-13, -1.269694e-14, 
    1.365391e-14, 3.515552e-13, 3.365082e-13, 4.364823e-13, 5.08276e-13, 
    8.147144e-14, -1.20879e-13, -4.525645e-14, -7.482133e-14, -5.15647e-14, 
    -4.714882e-14, -3.551565e-13, -4.378567e-13, 1.129953e-13, -2.916214e-13, 
    -4.834137e-13, -5.756528e-13, -3.45207e-13, -3.659763e-13, -2.535292e-13, 
    3.379495e-14, 1.448639e-15, 1.156343e-13, -6.639112e-14, -1.475373e-13, 
    -7.777074e-14, 1.597339e-13, 1.75372e-13, -1.632177e-13, 1.229446e-13, 
    -1.424939e-12, -1.636474e-13, -7.481446e-15, -9.825094e-14, 2.751141e-13, 
    3.288426e-13, -1.475353e-12, -5.547576e-13, 6.003325e-13, 5.53324e-13, 
    -3.28755e-13, 6.571069e-14, 9.064621e-13, 1.65586e-12, -3.411139e-13, 
    -1.724678e-12, 6.976526e-13, -2.053206e-12, -8.332652e-13, 2.069915e-12, 
    4.263444e-13, -2.141845e-13, -7.046172e-14, -8.877225e-14, -8.168915e-14, 
    3.427659e-13, 3.711867e-13, 4.655333e-13, 1.06277e-14, 6.649047e-14, 
    1.040113e-12, -1.212617e-13, 1.16238e-13, -1.312619e-13, 3.504324e-13, 
    -1.917098e-12, 2.726244e-13, 1.163058e-12, 5.357445e-12, -1.255167e-12, 
    -6.589441e-13, -6.300182e-13, 2.03676e-12, -4.352792e-13, -7.649813e-14, 
    -8.416533e-14, 1.048197e-12, 1.236141e-13, -1.362521e-13, 1.215567e-12, 
    -2.247082e-13, -4.10491e-13, 6.470719e-13, 1.065527e-13, 2.170069e-14, 
    2.357637e-13, -1.200364e-13, 4.927435e-13, 2.742473e-14, -1.380764e-12, 
    -8.554897e-13, 4.010703e-13, 1.082983e-12, -4.119054e-12, -2.587609e-13, 
    -2.860347e-13, -2.804603e-13, -1.819245e-12, -9.220458e-13, 1.0074e-13, 
    3.113817e-13, 4.4472e-13, 2.647234e-13, 1.172322e-15, 2.420348e-13, 
    -1.735081e-12, -5.309567e-12, 8.833608e-12, -3.888623e-15, 2.787427e-13,
  -4.46726e-14, -4.338196e-14, -2.569472e-14, -2.779027e-14, -1.348435e-13, 
    -2.481695e-13, -2.820313e-13, -8.719414e-14, 3.56451e-14, -1.079692e-14, 
    4.236889e-14, -5.827977e-14, -3.093706e-13, -1.630779e-13, 1.004058e-14, 
    1.18662e-14, -1.967801e-13, -2.429099e-13, -4.830129e-13, -3.098286e-13, 
    -4.512918e-13, -7.328235e-13, -4.975256e-13, -1.16164e-13, -2.864167e-13, 
    -4.893516e-13, -5.554654e-13, -1.060402e-13, -7.181755e-15, 5.30756e-14, 
    -8.437695e-15, -1.253234e-13, -2.140996e-13, -1.691702e-13, 4.862777e-14, 
    3.679695e-14, -8.035003e-13, 8.403868e-14, -3.587408e-14, -8.6363e-13, 
    1.446358e-12, -2.425005e-13, -5.909561e-13, -5.662701e-14, 4.415912e-14, 
    8.403694e-14, -1.083689e-12, -1.021117e-12, -1.324912e-14, 5.505735e-13, 
    -2.49167e-13, -1.131657e-12, -7.668658e-14, -2.05356e-11, 2.27568e-13, 
    -4.809625e-13, -4.029554e-13, -6.986744e-13, -8.274249e-13, 4.256213e-13, 
    -5.18488e-13, -1.230391e-12, -1.350864e-13, -1.13215e-13, -2.335618e-13, 
    1.510736e-13, -2.195466e-14, -3.891332e-14, 1.25025e-13, -4.557882e-13, 
    1.825227e-12, 2.966447e-13, -8.928969e-13, -1.381534e-13, 3.850725e-13, 
    -2.416692e-12, -5.253359e-13, 2.896555e-13, 9.549034e-12, -6.226963e-13, 
    6.946596e-13, 4.051416e-13, -1.05084e-12, 7.290696e-14, -2.254308e-13, 
    -5.380071e-13, -3.817155e-13, 4.738779e-13, -4.969379e-13, -1.677141e-12, 
    -2.795611e-13, -1.489961e-13, 5.193779e-13, -3.455562e-12, 4.239664e-15, 
    8.901248e-13, -2.702449e-13, 1.197584e-13, 1.019254e-13, 4.843491e-12, 
    -2.501888e-13, -5.586668e-13, 8.513164e-13, -2.156674e-12, 1.701278e-13, 
    1.008624e-12, 1.37753e-12, 2.572088e-12, 2.767002e-12, 2.116585e-12, 
    1.275216e-12, 8.284762e-13, 8.89934e-13, 6.521658e-13, 3.825551e-13, 
    1.059052e-12, -2.426478e-12, 1.737619e-11, -1.639422e-12, -7.907841e-13,
  -1.715017e-13, -1.781908e-13, -3.192169e-13, -4.317657e-13, -4.679451e-13, 
    -4.719558e-13, -3.518852e-13, -4.769796e-14, 1.127154e-13, 2.997325e-13, 
    1.67491e-13, 1.424971e-13, 4.571621e-13, 8.527484e-13, 6.028511e-13, 
    -7.677886e-14, -1.543599e-13, -3.95059e-13, -2.913746e-13, -7.4378e-13, 
    -3.383682e-13, 8.776313e-14, -5.335732e-13, -4.300588e-13, -1.024181e-13, 
    3.761574e-13, 3.913536e-15, -5.218881e-13, -3.773648e-13, -2.637057e-13, 
    4.74551e-13, 3.000239e-13, 4.956036e-13, -2.003814e-13, -1.609823e-14, 
    -2.430001e-14, -1.191162e-12, 7.098384e-13, 5.945661e-13, -7.507856e-13, 
    9.400952e-13, -6.142586e-13, -8.484324e-13, -1.534107e-13, 3.552714e-14, 
    8.409662e-13, -3.175724e-13, -8.959396e-13, -5.577844e-13, -1.040015e-12, 
    -1.258951e-12, -1.290384e-12, 3.34166e-13, -5.750275e-12, 5.877343e-13, 
    1.837912e-12, -1.033994e-11, 4.236112e-13, -9.545975e-14, 1.121856e-12, 
    -7.104317e-13, -7.99541e-13, -7.507883e-15, -2.883277e-13, -1.561667e-13, 
    -9.46937e-13, -1.106226e-12, -1.600525e-13, 1.161987e-13, -3.744366e-13, 
    4.636291e-13, -3.902434e-13, -7.252116e-13, -3.15456e-13, -3.137809e-13, 
    -1.01405e-13, -1.666306e-13, 1.473058e-12, -6.28713e-12, 5.426215e-15, 
    1.556047e-13, -1.787683e-12, -9.264811e-13, 8.352624e-13, 1.013495e-13, 
    -3.962386e-13, -3.211736e-13, -9.016399e-13, -4.517203e-13, 
    -5.071221e-13, -4.257011e-13, -4.824113e-13, 4.401271e-13, -7.403106e-14, 
    1.647849e-13, -5.497958e-12, -5.699968e-13, 2.685352e-13, -1.524308e-12, 
    -1.315828e-12, 1.010747e-12, -7.524155e-13, 5.252587e-13, 1.168805e-13, 
    2.999961e-13, 3.865103e-13, 5.5983e-13, 9.43412e-13, 6.038642e-13, 
    1.901534e-13, 6.307593e-13, 9.522938e-14, 1.064149e-13, 1.709743e-14, 
    -3.124445e-13, 2.990454e-12, 7.526833e-12, -5.433336e-13, -4.679859e-13, 
    -2.68327e-13,
  -1.490336e-13, -2.661898e-13, -1.681155e-13, -2.211148e-13, -2.184364e-13, 
    -2.563089e-13, -3.18634e-13, -1.965095e-13, 6.415007e-13, 1.037129e-12, 
    2.944173e-13, 1.073058e-12, 3.459594e-13, 1.175865e-13, -2.603334e-13, 
    -1.855169e-13, -5.337758e-13, -8.531023e-13, -4.812539e-13, 
    -7.746859e-13, -1.210726e-12, 2.435274e-13, -3.312489e-13, -1.57277e-13, 
    -7.101264e-14, -3.208545e-14, 5.538764e-13, -1.661588e-13, -3.013145e-13, 
    -1.414702e-13, -5.421913e-13, 9.885981e-13, -5.920264e-14, 7.145673e-13, 
    -1.438072e-12, -6.336043e-13, -6.148012e-13, -5.790247e-13, 3.955863e-13, 
    -7.225387e-13, -2.430195e-13, -4.149736e-13, -4.359048e-13, 
    -6.803681e-13, 1.965886e-12, 6.872281e-14, -6.717127e-13, -6.240251e-13, 
    -3.42551e-13, 1.517465e-11, 2.742025e-13, -1.904685e-12, -4.501524e-13, 
    -5.651535e-13, 5.88182e-13, 3.692296e-12, -1.253844e-12, -1.546804e-13, 
    -1.527833e-13, 2.073314e-12, -2.053913e-14, -4.703737e-13, -2.582934e-13, 
    -4.072825e-13, -5.401096e-13, -6.847439e-13, 1.517814e-13, -1.178224e-14, 
    -1.439265e-13, 2.085693e-13, 6.050022e-13, -2.842171e-14, -1.651776e-12, 
    -1.025638e-12, -8.928747e-13, -2.995659e-13, -4.347946e-13, 
    -4.167049e-13, -6.145405e-12, -8.344714e-14, 1.214528e-12, 3.031297e-13, 
    -6.052797e-14, -1.687983e-12, -4.597572e-13, 1.275008e-12, -1.30812e-13, 
    -6.24889e-13, -6.84155e-13, -6.694853e-13, -2.677025e-13, 3.145156e-12, 
    5.370045e-13, 1.145574e-12, -2.871731e-13, -8.748293e-13, -2.681077e-13, 
    -2.713108e-14, 2.702324e-12, -3.585049e-13, 1.999484e-12, -1.972502e-12, 
    6.757372e-13, 1.63783e-12, -5.095924e-13, 5.002804e-13, 8.642392e-13, 
    1.082606e-13, -5.203338e-13, -8.144735e-13, -4.736905e-13, -8.37358e-13, 
    -4.20039e-13, 2.695066e-14, -1.319334e-12, 2.299606e-12, -3.486642e-12, 
    -1.450584e-11, -2.259339e-12, -4.344303e-13,
  -5.014045e-14, -1.467021e-13, -2.051276e-13, -1.574157e-13, 7.659151e-14, 
    2.899486e-13, 8.693185e-13, -2.928213e-15, 1.43062e-12, 5.015294e-13, 
    3.579081e-14, 5.379169e-13, 3.118339e-14, -6.118023e-13, -7.369522e-13, 
    -1.375114e-12, -1.370326e-12, -5.080936e-13, -8.148066e-13, 
    -6.094708e-13, -4.766049e-13, 9.028195e-13, -9.083428e-13, -1.087033e-12, 
    -1.335446e-12, -4.106424e-12, -4.963821e-12, -3.620784e-12, 
    -2.749537e-12, -9.200557e-13, -1.839875e-12, 1.72394e-12, 1.894665e-12, 
    -1.010719e-13, -5.521555e-13, 5.599687e-14, 6.612766e-14, -5.897609e-13, 
    -8.229112e-13, 2.033929e-14, 7.28037e-13, -3.233289e-12, -6.614848e-13, 
    -1.535575e-12, 5.857106e-12, 2.761777e-12, 3.127776e-13, -4.784922e-13, 
    1.07708e-12, 2.968486e-11, 1.17175e-12, -2.614672e-12, 1.537548e-13, 
    -6.149112e-12, 5.117032e-13, 1.718903e-12, 3.448491e-13, -9.467454e-13, 
    4.826695e-15, 1.185156e-12, 1.367309e-12, -1.241091e-13, 1.604342e-12, 
    -6.885464e-13, -5.19021e-13, -5.849904e-13, -7.237266e-14, -1.254316e-12, 
    1.670844e-12, 2.431763e-12, 3.554518e-13, 2.961201e-12, -2.207665e-12, 
    -6.126072e-13, -1.789599e-12, 1.131456e-13, -4.699227e-13, -8.101367e-13, 
    2.628998e-12, 1.072073e-12, 1.946152e-12, 1.203538e-12, 5.793976e-14, 
    -1.642145e-12, 1.219649e-12, -5.308948e-13, 7.241444e-12, 1.408595e-14, 
    -8.604922e-14, 5.291184e-13, -4.292539e-13, 1.598779e-12, -2.275263e-14, 
    2.138706e-13, 2.120956e-12, -5.203332e-12, -1.318998e-12, -2.550876e-13, 
    2.805887e-11, 8.588047e-13, 5.31207e-12, 1.614996e-12, 1.571814e-12, 
    1.501826e-12, -5.992845e-13, -4.720807e-13, -8.526652e-13, -1.650444e-12, 
    -1.449382e-12, -1.353903e-12, -9.916096e-13, -1.166303e-12, 8.595208e-13, 
    4.179851e-13, -1.751863e-12, 1.999934e-12, -2.44392e-12, -1.083535e-11, 
    -1.065681e-12, -2.377029e-12,
  5.953293e-13, 6.129819e-13, 7.261136e-13, 9.378331e-13, 4.843348e-14, 
    -9.588441e-13, 7.374656e-13, 1.450645e-12, 1.062789e-12, 1.710798e-12, 
    1.431411e-12, 2.63406e-12, 4.596074e-12, 3.817419e-12, -4.752393e-12, 
    -2.198094e-12, -5.45447e-13, -2.318673e-12, -1.69403e-12, 1.290357e-13, 
    4.970191e-13, -6.896983e-13, -2.266992e-12, -9.938161e-13, -6.554091e-12, 
    -6.465134e-12, -8.093887e-12, -1.455525e-11, -7.014112e-13, -4.55147e-12, 
    -8.836099e-12, -3.972822e-12, 4.684114e-12, -5.042161e-12, 4.445611e-13, 
    2.682049e-12, -6.049799e-13, -5.627859e-13, 1.088851e-13, 1.480233e-13, 
    -4.15018e-13, -8.977902e-12, -2.462822e-13, -3.895914e-12, -1.797229e-12, 
    2.264661e-12, 6.841055e-13, -6.488837e-13, 8.917644e-13, -1.692958e-12, 
    1.335571e-12, 5.098422e-13, -6.272121e-13, -1.071476e-13, -7.614041e-13, 
    -3.421985e-13, 7.117085e-13, 1.049272e-13, 5.282996e-13, 3.815285e-12, 
    -2.214839e-12, 2.015554e-12, 5.803746e-12, -3.409328e-13, -5.16287e-13, 
    4.95104e-12, -2.751466e-12, 1.243808e-11, -4.060363e-13, -2.695649e-12, 
    -2.244399e-12, 1.157191e-11, -2.122053e-12, 1.053047e-13, -1.513761e-13, 
    4.695966e-13, -2.108383e-14, -2.813069e-12, -2.201828e-12, 6.172313e-12, 
    -1.690703e-12, -1.862642e-13, 6.080136e-13, -3.849976e-13, -1.477374e-12, 
    2.946865e-12, 7.414014e-12, -7.263634e-14, 4.668006e-13, -1.534939e-12, 
    1.820988e-12, 1.629807e-14, -6.409456e-14, -3.675754e-13, -6.999401e-13, 
    -1.854575e-12, -1.514844e-13, 1.621758e-13, 9.611562e-12, 8.781309e-14, 
    7.00659e-12, 1.811053e-12, 5.069712e-13, -3.394125e-13, 3.616274e-13, 
    -2.076672e-13, -1.817158e-12, -2.926132e-12, -2.248229e-12, 
    -2.591427e-12, -1.884493e-12, -2.56653e-12, -4.494738e-12, -5.418804e-12, 
    -1.597311e-11, 5.748887e-12, 5.200403e-12, 7.294693e-12, -1.090985e-13, 
    9.141576e-13,
  1.065925e-12, -1.592892e-12, -2.456813e-12, -5.260403e-12, -9.084122e-12, 
    -1.248218e-11, -8.679391e-12, 2.444656e-12, 2.978029e-11, 2.191208e-11, 
    3.188289e-11, 2.364742e-11, 1.132389e-11, 1.431499e-11, -7.055911e-12, 
    5.145884e-13, -8.955426e-12, -6.644685e-14, 3.042358e-13, -1.041167e-12, 
    -1.45578e-12, -2.065736e-12, -1.219247e-12, -8.318346e-13, -8.449963e-12, 
    -1.678557e-11, -2.352435e-11, -9.261536e-12, 1.198625e-11, -4.496459e-12, 
    -1.417738e-11, 9.853229e-12, 1.109668e-12, -5.721867e-12, -2.833456e-12, 
    -4.139467e-13, 1.829859e-12, -6.123782e-13, 7.183049e-11, -4.611645e-13, 
    -4.736878e-12, -4.003908e-12, 1.184788e-12, 6.355947e-12, -4.941048e-13, 
    -2.483513e-12, -1.207312e-12, 2.014638e-13, -1.121125e-12, -6.063396e-12, 
    -3.301942e-13, 5.375145e-13, 1.124767e-13, 1.108711e-11, -4.838445e-12, 
    7.668866e-14, 1.00287e-11, -1.706191e-13, 4.949153e-13, -4.562219e-12, 
    -1.077194e-12, 7.015499e-12, 1.383227e-12, -6.599266e-12, -6.011292e-12, 
    1.390588e-11, 4.312606e-12, 1.360645e-11, 7.239764e-13, -1.407369e-11, 
    -4.56496e-12, 7.667256e-12, 2.084777e-12, -5.693779e-13, 8.966161e-14, 
    1.901812e-13, 9.956619e-14, -3.462924e-13, -2.412738e-12, -1.739386e-12, 
    -3.639281e-11, 1.092224e-11, -2.356754e-12, -2.5833e-11, -1.535438e-13, 
    8.960055e-12, 1.70447e-12, -3.153144e-12, -1.026919e-12, 2.384759e-13, 
    2.435274e-13, -5.001665e-13, 2.476214e-13, 1.919281e-12, -4.251044e-13, 
    1.923312e-12, -2.493317e-12, 6.790679e-13, -3.339384e-12, 5.103918e-13, 
    6.161627e-12, 5.978273e-13, -5.371988e-13, -3.127835e-12, -4.015566e-12, 
    -9.065526e-13, -1.427802e-12, -6.233625e-12, -1.019557e-11, 
    -8.426038e-13, -1.018896e-11, -1.346229e-11, -1.3263e-11, -1.076766e-11, 
    -1.400041e-11, 1.469316e-11, 7.764553e-12, -2.588693e-12, 9.711329e-14, 
    1.334383e-11,
  -1.542033e-11, -1.780515e-11, -5.5142e-12, -5.054568e-12, -8.738399e-12, 
    -3.749334e-12, 6.725415e-11, 7.477408e-12, -2.347089e-11, -2.886541e-11, 
    -5.205025e-11, 6.250556e-14, -5.079548e-12, 1.626532e-12, -2.380707e-12, 
    -5.320766e-12, -4.729211e-12, -8.824885e-13, -9.574008e-13, 4.513445e-12, 
    4.634737e-12, 4.638345e-12, 5.052292e-12, 1.442846e-11, -8.893608e-12, 
    1.511435e-11, -7.001622e-12, -2.354272e-11, -3.85042e-12, -3.043904e-11, 
    -1.967498e-11, 1.383721e-11, 5.954182e-12, -2.33924e-13, -1.567635e-12, 
    1.320438e-11, 2.572775e-12, -4.952497e-13, -7.574608e-12, -3.315681e-14, 
    2.80248e-12, -3.002043e-12, 2.631395e-12, 5.022154e-12, -1.439293e-11, 
    1.819989e-11, -1.66156e-12, -9.101886e-13, 9.263734e-12, 9.741399e-12, 
    -1.277617e-12, -4.092338e-12, -3.36825e-13, 8.519241e-12, -5.721597e-12, 
    6.661338e-15, -6.270262e-12, 4.128364e-14, 6.611877e-13, -1.147459e-11, 
    6.4318e-12, 6.184109e-12, -1.885436e-12, -3.496603e-12, -1.114275e-12, 
    4.897194e-13, 9.432899e-12, 6.89232e-12, 1.854356e-11, -3.527678e-12, 
    -8.231194e-13, -3.642198e-11, 2.747524e-12, -3.626266e-12, 6.922241e-14, 
    6.467049e-14, -1.254552e-13, -2.47454e-11, -3.86874e-12, 2.568556e-12, 
    -4.357764e-11, 7.697554e-12, -1.690703e-12, -1.182598e-11, -5.994649e-13, 
    5.290768e-12, -7.407408e-13, -1.251144e-11, 1.721227e-13, 4.422573e-13, 
    5.378031e-12, 2.041201e-12, 7.553819e-13, 2.224398e-12, -1.317069e-11, 
    -1.561917e-13, -2.827294e-12, -1.203487e-11, -8.15692e-12, -2.987277e-13, 
    -7.56073e-12, -6.783886e-12, 3.299791e-13, -1.154204e-11, -3.022693e-12, 
    1.639522e-12, 2.041201e-12, -1.069533e-12, -1.539746e-11, 1.76259e-12, 
    -2.640893e-11, -1.055139e-11, -3.522238e-12, 8.267942e-12, 2.707001e-12, 
    1.80541e-11, 4.274997e-12, -9.159253e-13, 3.943026e-14, 7.822465e-12,
  1.849554e-11, 2.794726e-11, 9.567347e-12, 6.716849e-15, -2.237666e-11, 
    2.752976e-11, 2.236356e-11, -1.09564e-11, -4.732609e-11, -2.410883e-11, 
    2.530182e-11, -9.118151e-12, 5.934697e-13, 4.570622e-12, 3.752665e-12, 
    -9.322587e-12, -3.52427e-12, 4.651945e-12, 3.105495e-12, 4.90763e-12, 
    3.947398e-12, 5.974554e-12, 9.965084e-12, 2.453593e-13, 8.290368e-12, 
    -3.991418e-12, -2.89635e-12, -8.982481e-12, 3.492928e-12, 2.086498e-12, 
    -3.214823e-11, -3.363726e-11, -1.205991e-11, -6.078305e-12, 3.803957e-12, 
    -7.198347e-11, -6.049605e-13, -4.238762e-13, -5.044271e-11, 
    -1.510497e-12, 1.479883e-12, -5.910605e-12, 4.783937e-12, -1.113726e-12, 
    5.162926e-12, 7.888412e-12, 1.818462e-12, -7.656514e-13, 2.342149e-12, 
    8.621836e-12, -1.35908e-12, -9.6399e-12, -2.504774e-12, 5.036194e-13, 
    -5.091613e-12, 4.544143e-13, -8.070489e-12, 9.113988e-13, 1.070288e-12, 
    -5.374791e-12, 2.514489e-12, -9.819923e-14, 2.358891e-12, -4.231982e-12, 
    -1.266098e-13, -6.193546e-12, -1.798112e-11, 1.377748e-11, 6.73317e-12, 
    -3.37777e-11, -1.274275e-11, -1.505307e-11, 7.809309e-13, 1.434702e-11, 
    3.169842e-12, 9.037215e-14, -1.060749e-13, -2.26678e-11, -3.701133e-12, 
    5.946466e-12, -3.445386e-11, 9.012361e-13, 4.005685e-13, -1.267758e-11, 
    -1.967887e-11, -4.688583e-12, -1.789846e-12, -1.847544e-11, 7.031233e-13, 
    8.731904e-14, 5.342282e-12, -1.747935e-12, 1.795022e-12, -2.088113e-12, 
    -1.077938e-11, 5.997352e-12, -5.85243e-13, -5.35727e-12, 1.513512e-12, 
    -1.592149e-12, -5.587808e-12, -4.519503e-12, 1.671715e-12, -9.987716e-12, 
    -2.627676e-12, 3.766487e-12, 1.329159e-12, 9.75825e-12, -4.670764e-12, 
    1.710521e-12, -2.067163e-11, 7.008283e-13, 2.234202e-11, 1.009426e-11, 
    -8.055223e-13, 3.715023e-12, 1.036032e-12, -9.996396e-13, 4.844521e-12, 
    -7.087664e-13,
  1.969308e-10, 2.940975e-11, -3.205775e-11, -4.567374e-11, -4.123923e-12, 
    8.563039e-12, -2.020628e-11, -4.669209e-12, 6.111223e-12, 3.031925e-11, 
    6.194378e-12, -3.531536e-11, -1.231609e-11, -1.550821e-11, -2.286504e-12, 
    -4.454726e-12, -3.212069e-12, 3.772066e-12, 1.006622e-11, 6.695533e-12, 
    6.984691e-12, 9.92556e-12, 1.324191e-11, 4.678369e-12, 2.339351e-12, 
    -5.916045e-12, 2.979506e-12, -1.7919e-12, 3.971712e-12, 9.505119e-12, 
    -2.97885e-11, -1.607752e-10, -2.404926e-11, -1.030254e-11, -4.930112e-12, 
    9.895029e-12, -1.009975e-12, -3.312489e-13, -8.207557e-11, -1.744033e-12, 
    -4.409251e-13, -1.659595e-11, 4.53948e-12, -1.007889e-12, 5.82201e-13, 
    -6.244172e-12, 1.313366e-12, 1.090739e-12, 4.461875e-13, 1.676995e-12, 
    -1.622223e-12, 3.008083e-11, -3.669731e-12, 3.804512e-13, -3.499391e-12, 
    3.581024e-13, -1.562112e-11, 1.641615e-12, -2.278788e-13, -3.655957e-12, 
    -9.276968e-12, 1.978973e-12, 2.468581e-13, -2.68271e-12, 4.536338e-12, 
    -1.54815e-12, -5.030165e-11, 7.904233e-13, -1.297651e-11, -5.680206e-11, 
    4.448719e-12, -9.533285e-11, 3.612943e-12, -4.689027e-13, 1.005714e-11, 
    -1.34337e-14, -1.375566e-13, 2.807769e-11, -1.194159e-12, -1.24678e-13, 
    -2.432243e-11, 2.628857e-12, 4.978934e-12, -1.113348e-11, -2.154998e-12, 
    1.340211e-11, -4.381828e-12, -1.101252e-11, -1.336943e-13, 1.874612e-13, 
    7.109424e-12, 5.173706e-12, 1.077138e-12, 2.597877e-12, 6.922407e-12, 
    1.214667e-11, -4.546141e-13, -5.053069e-12, 6.496637e-12, -2.658185e-12, 
    4.879208e-12, 9.306944e-12, 1.888368e-12, -3.872316e-12, 1.753436e-11, 
    2.294576e-11, 2.578276e-11, 2.070305e-11, -9.287571e-13, -4.664047e-12, 
    2.398193e-12, 1.595768e-11, 1.864742e-11, 1.606715e-12, -8.787082e-12, 
    -8.412548e-13, 2.635114e-13, -1.818212e-12, 6.102549e-12, -7.789658e-12,
  1.694711e-10, -4.595879e-12, -5.922673e-11, -2.817702e-11, -1.455147e-11, 
    -3.979572e-11, -5.881173e-11, -4.30499e-11, -6.421785e-11, -5.851708e-11, 
    8.569034e-12, -7.326917e-11, -3.588907e-12, -3.319167e-11, -2.456191e-11, 
    -4.542555e-12, -6.598555e-12, 1.077366e-11, 7.889203e-12, 3.024581e-12, 
    4.057199e-12, 1.141909e-11, 1.195288e-11, 1.916289e-11, 7.122691e-11, 
    -2.094191e-11, -5.726974e-12, 7.281509e-12, 3.679756e-11, -1.198575e-11, 
    3.255229e-11, -5.108921e-10, -8.300238e-11, 1.937706e-11, 2.807155e-11, 
    -8.223866e-12, 4.563905e-13, -2.467193e-13, 1.214728e-11, 1.246614e-12, 
    -9.137135e-14, -2.640321e-11, 1.088934e-12, 3.211927e-13, -3.199008e-11, 
    -1.938194e-11, 3.868017e-13, -2.14273e-13, 3.492762e-13, 2.498002e-14, 
    -7.903164e-12, -2.554179e-12, 4.698686e-13, 1.145595e-12, -1.752484e-12, 
    2.416956e-13, 3.688239e-11, 1.257516e-12, 1.302128e-11, 6.049564e-12, 
    -1.325973e-11, -3.923528e-13, -2.584599e-13, -2.743583e-12, 1.091505e-12, 
    -1.378575e-11, -9.411805e-11, -3.993927e-11, 5.766165e-12, -1.130618e-11, 
    -2.825484e-11, 2.941003e-11, 2.556744e-11, -1.630918e-13, 1.43032e-11, 
    -8.337775e-14, -1.10606e-14, 3.123693e-11, 9.834355e-14, -2.996381e-12, 
    -1.792932e-11, 2.91219e-12, 5.809797e-13, 3.240963e-12, 1.666123e-11, 
    5.965151e-11, -4.544365e-12, -3.874678e-13, -1.204736e-12, -1.456613e-13, 
    2.850475e-11, 6.745005e-12, -4.543033e-13, -6.383194e-12, -1.056955e-11, 
    1.31151e-11, 1.073297e-12, -4.128253e-11, 1.061762e-11, -1.280598e-12, 
    -4.841683e-12, 5.139909e-12, 1.569106e-12, -2.940079e-13, 7.711265e-11, 
    4.343037e-11, 4.735023e-11, 2.885081e-11, -2.307377e-12, -4.419243e-12, 
    6.012746e-12, 3.555145e-11, 1.805267e-11, 1.060485e-12, -4.921397e-12, 
    -6.034284e-13, -1.218192e-13, -1.49027e-12, 2.630604e-12, -1.539102e-12,
  8.380407e-12, -5.116796e-12, -3.71021e-11, -4.586909e-11, -5.254219e-11, 
    -6.537171e-11, -5.329781e-11, -7.297052e-12, -4.166756e-11, 
    -1.065459e-11, -6.017942e-11, -1.864944e-10, 1.420686e-11, 3.74567e-12, 
    -1.418523e-10, -8.808065e-12, -6.657563e-12, 1.748046e-11, 6.925016e-12, 
    -7.850831e-12, -2.575495e-12, 1.338352e-11, 1.147682e-11, 2.224887e-11, 
    7.376899e-11, -1.609468e-11, -9.514833e-12, 3.319656e-11, 9.269274e-11, 
    -1.674216e-12, 1.519753e-10, 2.079137e-11, -2.18674e-10, -4.282463e-11, 
    1.398806e-10, -2.308678e-10, 6.125323e-13, 8.268386e-14, 6.927858e-11, 
    1.021427e-12, 5.733503e-12, -3.911693e-11, -1.696476e-12, 9.599196e-13, 
    -1.03566e-10, 5.886402e-13, -2.627232e-12, 1.980638e-13, 4.367173e-13, 
    1.600942e-13, -1.763395e-11, 5.259304e-11, 6.711076e-13, 1.737543e-12, 
    -7.775614e-13, 1.714184e-13, -5.641465e-11, 9.847678e-14, 2.215286e-11, 
    1.542616e-11, 7.952528e-12, -4.160006e-12, 1.906475e-12, 2.743006e-12, 
    1.783653e-11, -1.109255e-10, -5.839884e-11, -1.205853e-10, -2.752465e-12, 
    3.921752e-12, -7.144529e-11, -1.532068e-10, -1.251088e-11, -8.738965e-11, 
    1.463341e-12, -1.714184e-13, 1.814382e-13, 1.939793e-11, 4.266421e-13, 
    -2.225997e-12, -1.525036e-11, -4.04532e-12, -4.905409e-12, -6.552647e-11, 
    2.426281e-12, 1.022427e-10, 7.515388e-11, 4.474421e-12, -1.167975e-12, 
    -3.438361e-13, 6.408385e-11, 6.663026e-12, -1.168676e-12, -6.301692e-12, 
    -2.904299e-11, 1.047666e-11, 1.354028e-13, -9.496492e-11, 1.919442e-11, 
    1.695977e-13, -5.323564e-11, 5.073816e-12, 1.224507e-12, 1.949135e-13, 
    1.820513e-10, 8.664847e-11, 6.140977e-11, 3.313838e-11, -1.106271e-11, 
    -1.582268e-11, 6.074252e-12, 4.393441e-11, 2.742162e-11, 3.573364e-12, 
    8.026468e-12, 1.32272e-13, -6.900036e-14, -3.804665e-13, 5.741935e-13, 
    1.842815e-11,
  -3.54119e-11, -2.42697e-11, -5.27669e-11, -8.178369e-11, -9.56184e-11, 
    -7.480838e-11, -4.704259e-11, 2.328338e-11, 3.016987e-11, -9.354539e-11, 
    -1.381906e-10, -1.583509e-10, 8.536261e-11, 5.853074e-11, -1.943572e-10, 
    -9.833645e-12, 3.96887e-12, 1.786304e-11, 8.140877e-12, -2.312661e-11, 
    -3.465006e-12, 7.242429e-12, 1.87026e-11, 6.732592e-11, -8.013123e-11, 
    -6.746137e-11, -1.37701e-11, 3.345657e-11, 1.227056e-10, 5.000556e-11, 
    2.256775e-10, -1.184415e-10, 6.146572e-11, 1.183609e-11, 2.827671e-11, 
    1.357026e-11, -1.068701e-12, 2.832179e-13, -5.225376e-12, 5.970335e-13, 
    -1.223808e-11, -4.086265e-11, -8.836043e-12, 6.140435e-13, -2.428557e-10, 
    1.309952e-11, -6.92868e-12, 3.606559e-12, 5.550671e-13, 2.754186e-13, 
    1.125067e-11, 9.049894e-11, -6.933121e-13, 2.998801e-12, -7.617351e-13, 
    2.242651e-14, 3.262501e-12, -5.057732e-13, -5.449507e-12, 1.570849e-11, 
    4.078538e-11, -3.787703e-11, -1.22331e-11, 2.690821e-11, 3.033631e-11, 
    -1.445917e-10, -2.258038e-11, -2.223641e-10, -3.325851e-11, 3.987899e-11, 
    2.145173e-12, -3.70495e-10, -2.470986e-10, 1.722844e-12, -8.181057e-12, 
    -5.158096e-13, 9.525714e-14, 1.933309e-11, 4.105827e-13, -2.524891e-11, 
    -1.419553e-11, -1.385744e-11, -6.427747e-12, -1.841547e-10, 
    -3.389089e-11, -4.66166e-10, -1.359111e-10, 3.512524e-12, -4.770975e-13, 
    1.776357e-14, 7.276246e-11, 2.534906e-12, -6.702416e-13, 1.496581e-12, 
    -4.807199e-11, 5.297762e-12, -4.193668e-12, 4.7091e-11, 2.814748e-11, 
    2.239497e-12, -1.142613e-10, 8.234882e-11, 5.870582e-13, 1.637857e-13, 
    2.825116e-10, 2.521199e-10, 1.283784e-10, 6.247425e-11, -1.615841e-11, 
    -3.01219e-11, 1.629585e-12, 4.646616e-11, 3.083866e-11, -3.951728e-12, 
    1.347256e-11, 5.053735e-14, 2.384759e-13, 7.294165e-14, 2.602918e-13, 
    1.369771e-11,
  -5.745782e-11, -3.415379e-11, -8.151591e-11, -1.133722e-10, -1.160829e-10, 
    -8.997314e-11, -5.028844e-11, 1.571847e-10, 2.306157e-10, -3.010052e-10, 
    -2.34248e-10, -9.222378e-11, 1.585125e-10, 1.611469e-10, 1.400879e-12, 
    -6.224132e-12, 1.277862e-11, 4.176282e-11, -1.053957e-11, -3.150613e-11, 
    -6.382228e-12, 5.680123e-12, 2.56517e-11, 2.954303e-12, -9.87288e-11, 
    2.611444e-11, -2.078226e-11, 1.143807e-10, 2.377798e-10, 3.021452e-10, 
    2.926044e-10, 4.700174e-11, -1.710585e-10, -1.203293e-10, -3.291478e-11, 
    1.839855e-10, -3.34448e-12, 3.455014e-13, -5.082652e-10, 7.08722e-13, 
    -4.062666e-11, -1.338285e-11, -1.14575e-11, 6.339373e-13, -2.500433e-10, 
    1.095057e-11, -1.2496e-11, 3.081979e-12, 3.792966e-13, 5.094813e-13, 
    4.690881e-11, 5.654521e-11, 8.653921e-12, 5.164269e-12, 1.695755e-13, 
    -9.614531e-14, -1.05892e-10, -4.320544e-13, -3.455738e-11, 8.774093e-12, 
    6.476708e-11, -1.472358e-10, -1.554319e-10, 2.787801e-11, 2.19377e-11, 
    -1.537541e-10, -1.967737e-11, -4.277367e-10, -1.221101e-10, 1.203608e-10, 
    2.476004e-10, -4.045659e-10, 2.115439e-10, 3.55691e-11, -1.818275e-11, 
    -7.183143e-13, -4.818368e-14, 1.1531e-11, 2.023337e-12, -1.006615e-10, 
    -1.45286e-11, -9.839529e-12, -2.515543e-12, -1.9227e-10, -1.443048e-10, 
    -3.306162e-10, 1.544476e-11, 4.827472e-12, -1.849493e-13, -5.926371e-13, 
    1.241809e-10, 1.786558e-11, -6.328271e-13, 1.214224e-11, -7.164913e-11, 
    -3.133538e-12, -1.077232e-11, 1.37325e-10, 3.432743e-11, 4.440581e-12, 
    -2.088174e-11, 1.213241e-11, 2.68674e-13, 2.264855e-13, 3.09065e-10, 
    4.430138e-10, 3.133789e-10, 1.337936e-10, -1.959566e-11, -3.4867e-11, 
    9.170442e-14, 3.658962e-11, 2.136002e-11, -9.852341e-12, 8.406831e-12, 
    -2.294609e-13, 3.500533e-13, -1.439959e-13, -4.892753e-13, -7.427281e-11,
  -2.723288e-11, -4.596279e-11, -1.230238e-10, -1.273173e-10, -1.070526e-10, 
    -1.135336e-10, -2.055112e-11, 2.452292e-10, 5.653278e-10, -2.279701e-10, 
    -3.154992e-10, 3.758993e-11, 1.896736e-10, 2.621809e-10, 3.574918e-13, 
    -3.129052e-13, 1.073319e-11, 7.519585e-11, -4.115142e-11, -2.743894e-11, 
    -6.300294e-12, 1.031397e-11, 3.118084e-11, -1.456519e-10, 2.706724e-12, 
    -1.396594e-10, 5.882095e-11, 1.938747e-10, 6.26565e-10, 5.132184e-10, 
    5.693317e-10, 3.980238e-11, -5.81184e-11, -2.35659e-10, 1.484382e-10, 
    3.912324e-10, -5.171419e-12, 3.280709e-13, -5.753784e-10, -5.918643e-12, 
    -8.406689e-11, 1.602585e-11, -4.502843e-12, 2.413417e-12, -1.146501e-10, 
    1.270406e-11, -2.229816e-11, -2.470202e-11, 1.316014e-12, 6.574186e-13, 
    -1.073241e-11, -7.044099e-11, 2.016778e-11, 9.972201e-12, 1.887801e-12, 
    1.221245e-13, -2.225886e-10, 1.424194e-12, -6.004299e-11, 3.85133e-11, 
    6.859802e-11, -2.164096e-10, -3.910068e-10, 2.04845e-11, 3.403509e-11, 
    -1.372014e-11, -1.520912e-10, -6.806391e-10, -2.36303e-10, 8.200152e-11, 
    4.040683e-10, -5.366299e-10, 5.586509e-11, -8.333734e-11, -1.021041e-11, 
    -1.390443e-12, -3.341771e-14, -4.665379e-12, 3.595213e-12, -1.435079e-10, 
    -1.614175e-11, 4.567458e-12, 5.792256e-12, -1.693805e-10, -3.222289e-10, 
    -2.657221e-10, -1.020557e-10, 6.301182e-12, -5.904166e-13, -7.25553e-12, 
    5.74345e-11, 1.197736e-10, 4.665157e-13, 2.431122e-11, -1.119593e-11, 
    -1.279439e-11, -1.548512e-11, 3.086553e-11, 3.589973e-11, 3.321521e-12, 
    1.53221e-10, -1.554418e-10, 2.856604e-13, 7.180367e-13, 3.218648e-10, 
    3.813763e-10, 6.223808e-10, 2.950808e-10, -5.921041e-12, -3.439515e-11, 
    2.642331e-13, 1.573186e-11, -3.811618e-12, -5.901502e-12, -3.679279e-12, 
    -2.398082e-14, -8.670842e-14, -7.264744e-13, -2.772782e-12, -3.135816e-10,
  1.30397e-10, -3.642775e-11, -1.765059e-10, -1.478533e-10, -1.434604e-10, 
    -1.716796e-10, 5.391243e-12, 2.244835e-10, 7.340049e-10, 9.542411e-11, 
    -4.11438e-10, 2.083151e-10, 1.600693e-10, 3.183107e-10, -4.131628e-11, 
    1.025082e-11, 6.092549e-12, 9.670842e-11, -5.025602e-11, -1.475797e-11, 
    3.224088e-12, 1.288747e-11, 1.907274e-11, -1.84647e-10, -3.379164e-11, 
    -5.494218e-10, 4.636274e-10, 7.469225e-11, 1.103e-09, 7.605561e-10, 
    1.292459e-09, -5.633005e-11, 7.885248e-11, -6.307932e-10, 5.753797e-10, 
    3.246932e-10, -3.365663e-12, 6.348255e-13, -7.636611e-10, -2.861675e-11, 
    -8.695373e-11, 1.77085e-11, 8.779644e-12, 4.768158e-12, -1.48022e-10, 
    3.246114e-11, -2.986766e-11, -2.733103e-11, 3.22089e-12, 5.193623e-13, 
    3.979372e-11, -3.90914e-10, -3.332445e-13, 2.117808e-11, 1.073586e-12, 
    1.811884e-13, -1.676579e-10, 2.676259e-12, -1.26572e-10, 1.534373e-11, 
    5.902479e-11, -6.160761e-11, -2.609664e-10, 3.084964e-11, 5.429932e-11, 
    1.17657e-10, -3.96426e-10, -9.720171e-10, -4.675886e-10, 8.586554e-11, 
    4.561507e-10, -1.406045e-09, 2.843592e-11, -1.403926e-10, 3.284928e-11, 
    -3.351985e-12, 2.68896e-13, -2.520339e-11, 2.208767e-12, -1.413536e-10, 
    -2.078249e-11, -4.883161e-12, 1.84901e-11, -9.290524e-11, -5.462386e-10, 
    -3.750351e-10, -9.133672e-11, 1.518252e-11, -3.42204e-12, -2.361222e-11, 
    -4.02629e-11, 1.942855e-10, 6.97975e-12, 4.96641e-11, 4.39826e-11, 
    -9.92415e-12, -1.822862e-11, -1.439879e-10, 3.113954e-11, 1.577405e-13, 
    -1.534985e-10, -2.384802e-10, -7.361889e-13, 1.294964e-12, 2.821654e-10, 
    2.836131e-11, 6.599112e-10, 6.886918e-10, 2.058087e-11, -4.098055e-11, 
    1.076117e-11, -9.32765e-12, -1.882228e-11, 8.331114e-12, -6.050271e-12, 
    8.801848e-13, -1.121991e-12, -1.279088e-12, -5.218825e-12, -4.790923e-10,
  4.450236e-10, -1.88388e-10, -1.788703e-10, -1.684235e-10, -3.434515e-10, 
    -3.125002e-10, 7.140954e-13, 2.393623e-10, 5.802185e-10, -4.357901e-10, 
    -9.23448e-10, 1.908358e-10, 9.804424e-11, 3.138183e-10, 2.322409e-11, 
    2.68054e-11, -2.342659e-12, 1.111324e-10, -2.50715e-11, 7.633005e-12, 
    2.408207e-11, 1.670131e-11, 2.732037e-12, -8.291678e-11, -3.543779e-10, 
    -1.131427e-09, 2.685958e-10, 6.753016e-10, 1.620236e-09, 6.323262e-10, 
    2.122418e-09, 6.389076e-10, -2.073755e-10, 6.134666e-10, 1.534664e-09, 
    3.291891e-10, -9.78062e-13, 1.401768e-12, -2.094421e-09, -4.450147e-11, 
    -1.686828e-11, -1.021405e-11, 1.767431e-11, 7.903483e-12, -3.387264e-10, 
    6.52367e-11, -3.941114e-11, 1.067546e-11, -7.020873e-12, 5.218048e-14, 
    2.817757e-10, -8.331984e-10, -4.982628e-11, 3.443041e-11, -3.828582e-12, 
    7.904788e-14, -4.61494e-10, 2.334843e-12, -3.555737e-10, -3.255587e-10, 
    4.96545e-11, 2.078799e-10, 1.033573e-10, 3.950156e-11, 6.1004e-11, 
    7.428724e-11, -5.784493e-10, -6.705925e-10, -1.108793e-09, 1.568932e-10, 
    5.941239e-10, -4.003098e-09, -4.483152e-10, 1.624656e-11, 1.495549e-10, 
    -3.149481e-12, 8.437695e-13, -2.96918e-11, -2.606582e-12, -1.153833e-10, 
    -3.901324e-11, -2.468634e-11, 3.885336e-11, -3.298979e-10, -3.319514e-10, 
    -7.686118e-11, 1.138822e-10, 5.274536e-11, -1.218642e-11, -6.037659e-11, 
    -1.491216e-10, 2.287944e-10, 1.842126e-11, 6.563852e-11, -6.862599e-11, 
    5.404388e-12, -2.177671e-11, -2.556604e-10, 2.349054e-11, -1.163087e-11, 
    -8.36673e-10, -1.185146e-10, -3.718803e-12, -3.048006e-12, 2.529141e-10, 
    -1.232348e-10, 5.375043e-10, 1.198972e-09, 1.735323e-10, -4.777689e-11, 
    2.579448e-11, -2.789768e-11, -3.479528e-11, 1.551292e-11, 1.719869e-11, 
    2.458655e-12, 2.825296e-12, -1.785738e-12, -5.241474e-12, -2.939267e-10,
  5.397709e-10, 2.133156e-10, -1.37593e-10, -2.918874e-10, -6.741203e-10, 
    -6.387531e-10, -7.977263e-11, 2.587903e-10, 3.400729e-10, -1.974456e-10, 
    -5.920988e-10, 6.97149e-11, 6.273027e-11, 3.461373e-10, 2.313882e-11, 
    3.770211e-11, 4.625278e-12, 1.199396e-10, 1.405187e-11, 2.89937e-11, 
    5.559997e-11, 3.157652e-11, -4.554579e-12, -7.887024e-13, -8.898802e-10, 
    -1.915147e-09, -5.064145e-10, 2.323027e-09, 2.102428e-09, 2.215188e-10, 
    3.515879e-09, 1.422737e-09, -6.314238e-10, 1.263064e-09, 2.053532e-09, 
    4.281446e-10, 5.390177e-12, 1.897149e-12, -5.429406e-09, 3.426592e-12, 
    -1.556977e-10, -8.255796e-11, 1.401457e-11, 1.534955e-11, -2.686658e-09, 
    6.121681e-11, -7.229062e-11, 1.317533e-10, -3.378844e-11, 9.95648e-13, 
    3.963043e-10, -4.260592e-10, -1.415458e-10, 3.848655e-11, 1.699085e-13, 
    -5.506706e-14, -1.957311e-09, 2.08054e-11, -7.795393e-10, -2.324203e-10, 
    7.008083e-11, 3.030785e-10, 1.925677e-10, 3.017106e-11, 5.356995e-11, 
    -4.145555e-10, -4.33122e-10, -3.954916e-10, -1.316305e-09, -2.116458e-10, 
    6.505481e-10, -5.249408e-09, -6.043521e-11, 3.296314e-10, 5.201791e-10, 
    7.464251e-12, 1.957101e-12, -4.54925e-12, -1.079359e-11, -1.705018e-10, 
    -8.774848e-11, -6.198801e-11, 6.886403e-11, -4.793286e-10, -7.973355e-11, 
    5.615561e-10, 2.166587e-10, 1.076721e-10, -2.849815e-11, -1.418474e-10, 
    -3.733049e-10, 5.666145e-10, 2.850342e-11, 1.301725e-10, -3.803393e-10, 
    2.426255e-11, -2.631353e-11, -2.853362e-10, 1.580602e-11, -3.63336e-11, 
    -1.128946e-09, -4.124701e-11, -6.745715e-12, -1.685452e-11, 2.591314e-10, 
    3.041833e-11, 2.61263e-10, 1.48151e-09, -3.436895e-11, -9.153567e-11, 
    4.1954e-11, -5.124434e-11, -6.838619e-11, 4.785505e-12, 6.570033e-11, 
    3.798206e-12, 2.054579e-11, -1.232792e-12, -2.11009e-12, 3.208811e-11,
  5.276881e-10, 5.669101e-10, 5.892637e-10, 2.747989e-10, -4.369376e-10, 
    -1.007425e-09, -2.967901e-10, 2.438405e-10, 2.543139e-10, 2.127187e-10, 
    -3.645972e-10, -1.562732e-10, 2.386358e-11, 4.075567e-10, -4.217071e-12, 
    2.453788e-11, 2.768061e-11, 1.342748e-10, 4.217604e-11, 3.705125e-11, 
    8.199308e-11, 7.616663e-11, -1.776357e-14, 4.613199e-11, -1.447024e-09, 
    -2.684846e-09, -9.109762e-10, 2.39795e-09, 2.313133e-09, -3.197904e-10, 
    6.962164e-09, 2.43752e-09, -5.60977e-10, 2.030273e-09, 1.986759e-09, 
    1.165564e-09, -1.40119e-11, 4.385825e-12, -9.02352e-09, 9.05267e-11, 
    -2.719936e-10, -2.571845e-10, 7.620571e-13, 3.057798e-11, -2.323386e-09, 
    2.844658e-11, 8.972023e-11, 3.083045e-10, -5.839595e-11, 7.275069e-12, 
    2.190301e-10, 1.34342e-09, -1.46521e-10, 1.641709e-11, -1.582201e-11, 
    -4.618528e-13, -5.954472e-09, 9.387762e-11, -8.066557e-10, -1.434852e-10, 
    1.10699e-10, 2.075957e-10, -4.741914e-10, 1.219078e-11, 3.543121e-11, 
    -1.024585e-09, 4.944418e-10, 1.532747e-10, -1.619252e-09, 2.290541e-10, 
    -7.685586e-11, -4.047227e-09, -2.624283e-10, 1.089891e-09, 7.301885e-10, 
    3.207745e-11, 3.391065e-12, -4.837375e-11, -2.554099e-11, -2.490133e-10, 
    -1.801794e-10, -1.112667e-10, 9.580248e-11, -1.319076e-09, -4.233769e-11, 
    8.383942e-10, -1.342251e-10, 1.61922e-10, -5.359291e-11, -1.9973e-10, 
    -5.750955e-10, 1.427156e-09, 3.324097e-11, 3.23368e-10, -1.449234e-09, 
    2.680451e-11, -3.389644e-11, -8.145555e-10, 9.759304e-12, -4.109566e-11, 
    -8.34806e-10, 9.287149e-11, -7.499779e-12, -3.562928e-11, 3.69031e-10, 
    1.517471e-10, -2.48594e-10, 9.901058e-11, -2.068401e-09, -1.031179e-09, 
    5.743672e-11, -5.208634e-11, -1.725233e-10, -7.906564e-11, 1.761684e-10, 
    5.169909e-12, 6.324452e-11, 1.750378e-12, 9.41025e-13, 1.442864e-10,
  4.912302e-10, 5.681535e-10, 5.632508e-10, 7.643912e-10, 6.095782e-10, 
    -2.119087e-10, -3.015792e-10, 1.164473e-10, 5.966747e-10, -7.783996e-12, 
    -1.445979e-09, 3.706511e-10, -2.380318e-13, 3.227605e-10, -3.27784e-10, 
    -4.683684e-11, 4.997602e-11, 1.834017e-10, 5.820588e-11, 3.369749e-11, 
    8.143175e-11, 1.756639e-10, 6.039613e-14, 1.356035e-10, -1.289632e-09, 
    -3.364402e-09, -1.064404e-09, 3.393271e-09, 2.422286e-09, -1.255426e-09, 
    1.53858e-08, 4.946703e-09, 2.061746e-10, 2.704386e-09, 1.915243e-09, 
    6.278533e-10, -3.509584e-11, 8.583356e-12, 1.448885e-09, 4.791971e-11, 
    -1.03568e-10, -4.812186e-10, -2.786038e-11, 5.515211e-11, -3.633254e-10, 
    -1.4591e-11, 1.211138e-09, 3.875904e-10, -6.856667e-11, 3.19984e-11, 
    -2.531024e-10, 1.836856e-09, 3.391065e-11, -9.078675e-11, -7.918714e-11, 
    -1.552536e-12, -1.010691e-08, 2.159887e-10, 5.968204e-11, 6.586696e-10, 
    1.125251e-10, 6.359713e-11, 9.904007e-10, 1.715321e-11, 3.42915e-11, 
    -1.081386e-09, 3.163798e-10, -1.013767e-10, -4.711975e-09, -5.990408e-10, 
    -1.152966e-09, -1.672714e-09, 2.639418e-10, 3.111754e-09, 2.004426e-09, 
    6.035705e-11, 4.014566e-12, -1.459242e-10, -2.554898e-11, -1.642313e-10, 
    -3.132179e-10, -1.25944e-10, 8.931877e-11, -8.630547e-09, -6.498269e-11, 
    -2.119616e-09, -8.707666e-10, 1.990834e-10, -8.939982e-11, -4.229612e-10, 
    -6.816592e-11, 2.080444e-09, 3.13527e-11, 6.207834e-10, -2.530538e-09, 
    3.348788e-12, -5.377316e-11, -1.629044e-09, -6.419754e-12, -5.533636e-11, 
    2.133937e-10, 3.373586e-10, -3.553602e-12, -4.991829e-11, 4.378681e-09, 
    1.313687e-10, -2.79524e-10, 2.878018e-10, -2.103882e-10, -1.998512e-09, 
    3.179323e-11, -2.145484e-11, -4.056169e-10, -4.131202e-10, 3.097433e-10, 
    4.083489e-12, 9.899459e-11, 4.862777e-12, -4.987122e-12, 2.996003e-11,
  3.621459e-10, -7.507204e-10, 2.024176e-09, 8.892407e-10, 1.086615e-09, 
    8.412222e-10, 3.856506e-10, 1.369465e-10, 1.526413e-09, -1.971792e-10, 
    -2.22828e-09, 4.55729e-09, -4.576783e-10, 1.559997e-11, -9.83281e-10, 
    -5.559357e-11, 6.914647e-11, 2.315268e-10, 8.455103e-11, 2.456702e-11, 
    4.055423e-11, 3.137011e-10, 2.170708e-12, -3.656808e-11, -7.589769e-10, 
    -3.790422e-09, 1.306343e-09, 4.657121e-09, 3.391811e-10, -2.752873e-09, 
    1.38186e-08, 3.889706e-09, 2.006626e-09, 2.110166e-09, 1.513552e-09, 
    8.817658e-10, 1.670607e-10, 1.505285e-11, 3.917574e-09, -8.141988e-10, 
    3.685464e-10, -5.146212e-10, -1.202238e-11, 1.025362e-10, 1.482402e-09, 
    -2.166907e-10, 2.606459e-09, 4.124701e-10, -1.089354e-10, 4.774314e-11, 
    8.526158e-11, 2.738538e-10, -1.648953e-11, -2.501913e-10, -1.598078e-10, 
    -4.146017e-12, -1.546212e-08, 3.816943e-10, 9.221743e-10, -1.326761e-11, 
    5.556089e-11, -5.022471e-11, 4.380603e-10, 2.04345e-11, 7.6232e-11, 
    -2.444441e-09, -5.070468e-10, -8.157919e-10, -2.746408e-09, 
    -1.099924e-09, -1.588337e-09, -6.765539e-10, 2.954685e-10, 3.9723e-09, 
    4.476623e-09, 5.331557e-11, 2.303935e-12, -2.311005e-10, 2.117453e-11, 
    6.256293e-10, -4.583534e-10, -1.714998e-10, 1.174989e-10, -7.869534e-09, 
    -9.602026e-10, -8.18293e-10, -5.48031e-10, 1.956089e-10, -1.231311e-10, 
    -1.46709e-09, 8.971135e-10, 1.676522e-09, 3.09619e-11, 8.524118e-10, 
    -3.368502e-09, -3.146354e-11, -1.107288e-10, -2.469367e-09, 
    -3.177902e-11, -8.528574e-11, 4.134755e-10, 6.29174e-10, 6.087575e-12, 
    -6.291767e-11, 7.001102e-09, 1.423324e-10, 4.646594e-11, 1.274653e-09, 
    1.417131e-09, -6.650289e-10, -1.530971e-10, -2.784262e-11, -6.331824e-10, 
    -7.965077e-10, 4.270895e-10, 5.055512e-12, -7.409184e-12, -1.149747e-12, 
    -2.914824e-11, 2.499334e-11,
  1.142098e-09, -4.909111e-09, 6.014986e-09, 2.41279e-09, 4.074963e-10, 
    1.527809e-09, 9.101768e-10, 5.625509e-10, 2.847244e-09, 4.977494e-10, 
    -3.157709e-09, 3.304649e-09, 7.423608e-10, 1.072053e-09, -1.637176e-09, 
    -2.133163e-10, 1.712266e-11, 2.065761e-10, 1.355644e-10, -2.469847e-11, 
    -5.115908e-13, 4.562821e-10, -5.132961e-11, -2.089848e-10, -1.943718e-09, 
    -3.700563e-09, 1.175181e-09, 7.20199e-09, -2.929411e-09, -5.484551e-09, 
    4.531486e-09, 4.756387e-09, 5.775945e-09, 9.035261e-10, 5.172183e-10, 
    -7.482015e-11, 4.796504e-10, 3.392486e-11, 4.627267e-09, -2.35853e-09, 
    7.675879e-10, -9.859491e-11, 5.248424e-11, 1.252214e-10, 1.993072e-09, 
    -4.520189e-10, 4.401514e-09, 3.712941e-10, -3.030323e-10, 1.323652e-11, 
    6.957102e-11, 1.244871e-11, 4.013344e-10, -1.086875e-10, -2.58116e-10, 
    -7.851497e-12, -2.233584e-08, 6.71416e-10, 1.736392e-09, -6.265566e-10, 
    3.335288e-11, -2.118838e-10, -9.576695e-11, 3.701361e-11, 1.164466e-10, 
    -5.329781e-09, 6.361205e-10, -6.459317e-09, 1.433122e-09, -2.099384e-09, 
    -5.585434e-10, -2.476639e-09, 2.076632e-10, 2.768516e-09, 2.925923e-09, 
    9.947598e-14, 2.602363e-12, -3.171579e-10, -6.78211e-13, 2.01247e-09, 
    -5.894663e-10, -4.177426e-10, 2.854605e-10, -7.320978e-09, -1.147811e-10, 
    6.432828e-10, 6.040892e-10, 1.68626e-10, -4.616707e-11, -2.634877e-09, 
    7.09349e-10, 2.371812e-09, 4.076028e-11, 9.225559e-10, -4.177338e-09, 
    -7.901946e-11, -2.312618e-10, -3.047916e-09, -5.393019e-11, 
    -1.423871e-10, 5.582024e-10, 9.512826e-10, 9.838352e-12, -8.25997e-11, 
    6.718508e-09, 1.20906e-10, 1.022471e-10, -5.049401e-10, 8.495675e-10, 
    -5.345697e-10, -2.650609e-10, -9.677592e-12, -9.622028e-10, 
    -9.307115e-10, 5.442189e-10, 6.811262e-12, -4.024887e-10, -2.268541e-11, 
    -5.743583e-11, 7.247536e-12,
  3.27648e-09, 5.226493e-09, 3.081933e-09, -3.9444e-10, -1.792817e-09, 
    8.481855e-10, 2.011372e-09, 1.286619e-09, 3.289156e-09, 2.346891e-09, 
    2.831708e-09, -5.105143e-10, 2.250655e-09, 3.032707e-09, -2.192682e-09, 
    -7.56868e-10, -3.622496e-10, -3.97371e-11, -8.376944e-11, -1.11843e-10, 
    8.835599e-12, 4.099228e-10, -6.830092e-11, 1.385558e-13, -2.728317e-09, 
    -5.987921e-10, 1.632227e-09, 9.2767e-09, 4.375771e-10, -8.978478e-09, 
    6.557851e-09, 5.41527e-09, 6.473268e-09, -1.144887e-09, -4.530172e-10, 
    -2.308614e-09, 9.789595e-10, 4.958522e-11, 3.337785e-09, -1.208827e-09, 
    1.066646e-09, -8.359535e-12, -3.806768e-10, -7.239498e-11, -3.653646e-10, 
    -4.937171e-10, 8.678821e-09, 2.349374e-10, -7.710902e-10, -1.66823e-10, 
    7.934275e-11, -3.157687e-10, 8.31843e-10, -1.444178e-11, -3.229587e-10, 
    -8.842704e-12, -1.953905e-08, 1.633151e-09, 2.923243e-09, -4.769269e-10, 
    1.054126e-10, -4.662901e-10, -1.224727e-10, -9.98913e-10, 3.762111e-11, 
    -8.774126e-09, -6.878373e-10, -7.188053e-09, 6.386525e-09, -4.529799e-09, 
    6.046115e-10, -4.278181e-09, -1.416858e-10, 2.643954e-09, -3.063755e-10, 
    -5.960388e-11, 1.589839e-11, -3.828085e-10, -1.718874e-11, 2.652055e-09, 
    -6.745076e-10, -9.09273e-10, 5.969945e-10, -7.933981e-09, 2.007763e-09, 
    7.484822e-10, 2.282174e-09, 1.614602e-10, 3.153788e-10, -3.974865e-09, 
    -5.193819e-10, 2.770954e-09, 5.339373e-11, 8.863815e-10, -4.483386e-09, 
    -1.732481e-10, -3.850495e-10, -3.233797e-09, -1.029186e-10, 
    -2.189303e-10, -4.345146e-10, 1.130708e-09, -3.508305e-12, -1.017746e-10, 
    4.954497e-09, -4.3946e-10, 3.091678e-10, -9.808083e-10, -2.032753e-09, 
    4.135607e-10, 1.180521e-09, 9.062973e-12, -9.382326e-10, -5.065637e-10, 
    6.80668e-10, -1.734435e-12, -1.35099e-10, -5.116441e-11, -7.194245e-11, 
    -1.428226e-10,
  5.332595e-09, -5.899295e-09, -8.407852e-09, -3.003578e-09, -4.153804e-09, 
    -1.136044e-09, 2.636881e-09, 2.371792e-09, 3.125024e-09, 3.510905e-09, 
    8.441901e-09, 2.591264e-09, 2.963219e-09, 6.075908e-09, -2.642707e-09, 
    3.156316e-10, -5.824433e-10, -9.511467e-10, 6.209717e-10, -1.861338e-10, 
    2.728484e-11, 2.264073e-10, 1.961098e-11, -4.073115e-10, 3.558824e-09, 
    1.14386e-09, 2.042043e-09, 1.059703e-08, 2.844274e-09, -1.197134e-08, 
    1.076486e-08, 6.473243e-09, 1.138432e-09, -7.39476e-10, -6.218102e-10, 
    -3.872714e-09, 1.444519e-09, -4.561684e-12, 3.336737e-09, -6.898717e-10, 
    2.558647e-09, -4.01883e-10, -1.878526e-09, -9.972423e-11, 1.554326e-09, 
    3.871037e-11, 5.811117e-09, 3.117222e-10, -1.317318e-09, -2.176712e-10, 
    1.21851e-10, -2.063075e-09, 1.144807e-09, -1.788749e-10, -7.670479e-10, 
    -4.050094e-12, -2.27927e-08, 5.901015e-09, -1.293841e-09, 7.022862e-10, 
    2.24361e-10, -5.509548e-10, -5.665299e-10, -4.154583e-09, -6.737651e-11, 
    -1.429228e-08, 3.190451e-09, -3.950134e-09, 1.272181e-08, -7.505491e-09, 
    7.740084e-10, -3.295582e-09, -6.849632e-10, 3.038366e-09, 1.637429e-09, 
    -8.131451e-11, 3.695888e-11, -3.275389e-10, -4.694059e-11, 3.716622e-09, 
    -8.052154e-10, -1.349881e-09, 1.027431e-09, -1.050151e-08, -1.145594e-09, 
    5.334755e-11, 2.202938e-09, 2.115996e-10, 4.940151e-10, -5.801482e-09, 
    -2.281155e-09, 2.181838e-09, 5.333334e-11, 1.139267e-09, -8.141399e-10, 
    -2.484484e-10, -4.721414e-10, -1.063427e-09, -1.462865e-10, 
    -2.991953e-10, -7.710526e-10, 7.109584e-10, -5.469936e-11, -9.964829e-11, 
    3.24178e-09, -1.580617e-09, -2.505942e-10, -2.141434e-09, -5.837165e-09, 
    -1.441038e-09, 4.306372e-09, 1.675119e-09, -8.576535e-10, 8.441248e-11, 
    9.474661e-10, -4.059188e-11, -4.835243e-12, -4.577316e-11, -7.069367e-11, 
    -3.053628e-10,
  7.512028e-09, -1.70283e-09, -9.552451e-09, -3.633659e-09, -3.122437e-09, 
    -5.157489e-09, 2.629889e-09, 4.083091e-09, 2.470273e-09, 3.733561e-09, 
    1.180541e-08, 7.025108e-09, 4.954586e-09, 6.674128e-09, -3.200341e-09, 
    -8.663537e-10, -3.370133e-10, -2.095945e-09, 2.89133e-09, -2.158231e-09, 
    -4.587264e-11, -1.350031e-10, 5.857714e-11, -5.159393e-10, 1.475337e-08, 
    4.970275e-09, 2.044061e-09, 1.296277e-08, 6.799638e-09, -1.109487e-08, 
    1.821675e-08, 5.335494e-09, 7.45419e-09, -1.680178e-09, -6.452865e-10, 
    -5.266259e-09, 1.758647e-09, -1.335216e-10, 4.558245e-09, 2.323333e-10, 
    4.883833e-09, -6.159837e-10, -2.788767e-09, -2.354694e-11, -2.294769e-10, 
    4.796163e-10, -9.017896e-09, 1.454552e-10, -1.729035e-09, -1.645226e-10, 
    6.385648e-11, -4.726644e-09, 1.291238e-09, -1.832348e-10, -1.666948e-09, 
    -9.066525e-12, -2.904275e-08, 1.535949e-08, -1.518971e-08, 2.072177e-09, 
    2.553406e-10, -6.035634e-10, -1.115865e-09, -4.770015e-09, 3.840341e-11, 
    -2.065073e-08, 4.244384e-09, -1.858012e-09, 2.069527e-09, -7.95518e-09, 
    3.110756e-10, -1.690466e-09, -6.606911e-10, 1.715705e-09, 3.505068e-09, 
    -7.466383e-11, 5.070788e-11, -3.618013e-10, -7.393623e-11, 4.826916e-09, 
    -1.81609e-09, -1.32373e-09, 2.009699e-09, 3.473701e-09, 1.234156e-09, 
    1.716387e-10, 8.104166e-10, 3.446701e-10, -5.06005e-10, -9.086094e-09, 
    -6.554757e-09, 2.017686e-09, -5.82645e-13, 7.414573e-09, 1.875122e-09, 
    -2.744685e-11, -4.435265e-10, 2.094453e-09, -3.780087e-11, -3.668504e-10, 
    -3.692833e-10, -4.144773e-10, -1.216947e-10, -1.342997e-10, 
    -5.176105e-09, -1.350685e-09, -1.13701e-09, -4.568165e-09, -6.63556e-09, 
    -6.209802e-09, 8.75599e-09, 2.170992e-09, -1.049557e-09, 6.473613e-10, 
    1.850538e-09, -2.732463e-11, 2.789236e-11, 2.248335e-11, -6.837197e-11, 
    -4.103811e-10,
  8.162658e-09, -1.643912e-09, -4.8841e-09, -4.976698e-09, -1.469346e-09, 
    -6.926598e-09, 2.403624e-09, 5.868685e-09, 6.515393e-10, 3.263722e-09, 
    9.783832e-09, 1.22256e-08, 4.084654e-09, -5.534389e-09, 1.216961e-09, 
    -1.212669e-09, 3.265711e-10, -3.047489e-09, 6.310607e-09, -4.93327e-09, 
    -2.031584e-10, -4.560547e-10, -1.226681e-10, -4.276899e-10, 1.713477e-08, 
    1.300231e-08, 2.116053e-09, 1.036216e-08, 1.115762e-08, -1.099687e-08, 
    2.098506e-08, 5.313666e-09, 7.12015e-09, -1.789772e-09, 1.254534e-10, 
    -7.188646e-09, 1.495511e-09, -1.092957e-10, 8.327618e-09, 7.989467e-10, 
    7.325377e-09, -2.789875e-10, -1.68852e-09, 1.503766e-10, -1.284548e-09, 
    2.069612e-09, -2.486843e-09, 4.973799e-11, -2.95704e-09, -9.188028e-11, 
    -9.50493e-11, -3.704201e-09, 1.843529e-09, 5.079528e-11, -2.736097e-09, 
    -3.777245e-11, -3.258492e-08, 2.476975e-08, -2.183322e-08, 3.684832e-09, 
    3.719265e-10, -1.488104e-09, -1.759133e-09, -4.390984e-09, -1.535568e-10, 
    -1.563939e-08, 4.995002e-09, 6.487539e-10, -5.201173e-09, -9.150881e-09, 
    -2.474962e-10, -1.476735e-09, 1.620037e-10, -1.063995e-09, 1.762146e-09, 
    -1.658691e-10, 5.806555e-11, -3.760903e-10, 4.858697e-12, 7.317681e-09, 
    -5.315172e-09, -7.186955e-10, 3.715513e-09, 7.633957e-09, 2.552326e-09, 
    7.324843e-10, 9.764562e-10, 4.379217e-10, -2.69097e-09, -1.39089e-08, 
    -1.211998e-08, 2.637989e-09, -1.380727e-10, 1.889845e-08, -8.647589e-10, 
    6.393066e-10, -3.875812e-10, 4.671506e-09, 3.399236e-10, -4.108301e-10, 
    1.703825e-09, -1.112202e-09, -2.719425e-10, -2.485621e-10, -1.113335e-09, 
    -5.200036e-10, -1.445471e-09, -5.428603e-09, -5.924676e-09, 
    -4.412755e-10, 1.539894e-08, 8.363941e-10, -1.976389e-09, 1.275907e-09, 
    3.306127e-09, -7.997869e-12, 9.449508e-11, 1.171188e-10, -5.559286e-11, 
    -2.797833e-10,
  5.417007e-09, 7.015046e-10, -2.46331e-09, -3.939419e-09, -4.170033e-10, 
    -3.500702e-09, 1.491173e-09, 6.802054e-09, 4.268941e-10, 2.792945e-09, 
    6.156654e-09, 1.162329e-08, 1.952003e-09, -4.478977e-09, 2.1397e-09, 
    -1.431476e-09, 1.041923e-09, -3.753541e-09, 1.077343e-08, -2.641116e-09, 
    -1.791932e-09, -3.648779e-10, -1.043645e-10, -6.195933e-12, 7.112931e-09, 
    8.509062e-09, 3.556579e-09, 9.755013e-09, 1.37473e-08, -2.421558e-08, 
    2.421655e-08, 6.399034e-09, 1.413616e-08, -2.55335e-09, 2.950742e-10, 
    -1.039518e-08, 9.053736e-10, 1.151079e-10, 1.600051e-08, -5.345608e-10, 
    8.907875e-09, 2.540332e-10, -1.444917e-09, 3.576464e-10, 1.382602e-09, 
    1.136482e-08, 1.382253e-08, 1.816716e-10, -5.160541e-09, -3.760903e-11, 
    -4.943033e-10, -3.252467e-09, 3.2164e-09, 5.343295e-13, -3.306541e-09, 
    -4.553158e-11, -3.364943e-08, 3.23524e-08, -2.080411e-08, 3.762068e-09, 
    1.209344e-09, -2.591662e-09, -1.957915e-09, -6.757238e-09, -8.540383e-10, 
    2.623892e-09, 9.199255e-09, 4.974595e-09, -3.829371e-09, -1.281256e-08, 
    -1.028866e-10, -2.512877e-09, -1.209457e-09, -1.390731e-09, 3.453351e-09, 
    -2.262368e-10, 6.678391e-11, -7.090648e-10, 1.998004e-10, 1.130132e-08, 
    -1.131886e-08, -2.395779e-10, 5.775433e-09, 8.535039e-09, -1.399201e-09, 
    1.063256e-09, 2.071033e-09, 4.119443e-10, -3.521961e-09, -1.757343e-08, 
    -1.209776e-08, 4.968673e-09, -2.930705e-10, 1.542438e-08, -4.572371e-09, 
    1.051836e-09, -4.88376e-10, 7.904191e-09, 1.092872e-09, -4.614094e-10, 
    3.305615e-09, -2.255536e-09, -6.219985e-10, -3.368683e-10, 2.012484e-09, 
    3.921627e-10, -5.424567e-10, -2.757986e-09, -4.021899e-09, 3.095977e-09, 
    1.955306e-08, -7.661356e-10, -3.909975e-09, 2.151239e-09, 2.978538e-09, 
    3.012133e-11, 1.497966e-10, 2.112976e-10, -6.456347e-11, -6.252776e-12,
  3.465857e-09, 1.949331e-09, 9.770815e-10, 5.624656e-10, -1.213607e-10, 
    6.127152e-10, -3.69937e-10, 5.797631e-09, 2.116678e-09, -1.436433e-10, 
    4.822709e-09, 8.521226e-09, -4.06385e-09, 7.971039e-09, 6.643347e-09, 
    -1.010829e-09, 2.292569e-09, -6.747172e-09, 1.742308e-08, -1.524484e-09, 
    -5.615391e-09, -1.378453e-10, 2.852403e-10, 1.795684e-10, 1.07292e-09, 
    -3.57727e-09, 5.67502e-09, 3.103008e-08, 1.279852e-08, -4.52809e-08, 
    2.335508e-08, 8.550842e-09, 1.908853e-08, -3.547029e-09, -3.574655e-09, 
    -1.45705e-08, 1.104451e-09, 4.387317e-10, 2.16848e-08, -2.368756e-09, 
    9.148289e-09, 1.556145e-09, -2.04173e-09, 6.029346e-10, 8.355755e-09, 
    2.701199e-08, 3.129813e-08, 6.733814e-10, -7.868425e-09, -4.520828e-11, 
    -9.999681e-10, -3.617231e-09, 5.990802e-09, -1.696776e-10, -3.786222e-09, 
    9.379164e-12, -1.718359e-08, 3.830455e-08, -1.748519e-08, 2.59832e-09, 
    2.097636e-09, -3.047205e-09, -7.304379e-10, -6.886523e-09, -2.067486e-09, 
    -8.893721e-10, 2.68887e-08, 6.834057e-09, 1.0441e-09, -1.516753e-08, 
    4.970389e-10, -2.046136e-09, -1.581384e-09, -1.241915e-09, 7.471709e-09, 
    -2.662546e-10, 7.710099e-11, -2.024748e-09, 7.091501e-10, 1.286185e-08, 
    -1.598579e-08, -6.066515e-10, 7.394789e-09, 8.289419e-09, -3.838068e-09, 
    -1.663068e-09, 3.156913e-09, 2.447109e-10, -1.862094e-09, -1.672703e-08, 
    2.763898e-09, 8.471455e-09, -5.599787e-10, -1.379701e-08, -6.193659e-09, 
    -4.554238e-10, -7.772428e-10, 7.193023e-09, 2.151467e-09, -5.796096e-10, 
    2.862294e-09, -3.348354e-09, -9.60334e-10, -4.186909e-10, 6.937398e-09, 
    2.810111e-09, 1.883052e-09, -1.505725e-09, -5.69554e-09, 9.776329e-09, 
    1.737089e-08, -4.582148e-10, -7.638164e-09, 4.025537e-09, 1.169099e-09, 
    -1.127773e-11, 2.126939e-10, 2.150422e-10, -7.860024e-11, -2.131628e-11,
  1.064848e-09, 1.96826e-09, 1.27261e-09, 1.825242e-09, 6.565983e-10, 
    2.489514e-09, -5.931554e-09, 4.387459e-09, 3.159641e-09, -2.387651e-09, 
    2.732975e-09, 7.24441e-09, -1.242347e-08, 2.91169e-09, 8.761845e-09, 
    -4.436748e-09, 2.99587e-09, -1.001078e-08, 2.445363e-08, -3.754792e-09, 
    -8.034306e-09, -6.69047e-11, 6.48356e-10, -8.252528e-10, -6.28404e-10, 
    -2.080469e-09, 1.086806e-08, 3.29357e-08, 1.432994e-08, -4.612554e-08, 
    1.815437e-08, 1.148209e-08, 2.257832e-08, -2.961372e-09, -1.157179e-08, 
    -1.661141e-08, -8.46984e-10, 8.22439e-10, 2.399906e-08, -3.888104e-09, 
    7.673304e-09, 3.815046e-09, 3.583267e-09, 7.072281e-10, 1.077717e-08, 
    3.927192e-08, 4.565746e-08, 8.238317e-10, -1.1872e-08, -4.896705e-11, 
    -1.377067e-09, 3.896048e-10, 1.087675e-08, -4.02008e-10, -3.204236e-09, 
    1.338378e-10, -8.431584e-09, 4.214428e-08, -8.477656e-09, -2.886075e-09, 
    -1.191665e-09, -4.213973e-09, -1.637659e-10, -4.02938e-09, -3.339835e-09, 
    7.918857e-10, 1.405675e-08, -2.736499e-09, 2.143622e-09, -1.053257e-08, 
    8.155325e-10, 7.313076e-09, 2.042214e-09, -1.433534e-09, 1.417479e-08, 
    -2.248157e-10, 1.51708e-10, -3.612456e-09, 1.585846e-09, 8.413963e-10, 
    -1.712479e-08, -1.780636e-09, 8.218706e-09, 3.584944e-09, 1.955414e-11, 
    -3.780656e-09, 2.803517e-10, -3.211653e-11, 7.215153e-10, -1.373792e-08, 
    1.594077e-08, 1.173255e-08, -1.786034e-09, -3.50458e-08, -5.041954e-09, 
    -4.120449e-09, -1.199953e-09, -5.262564e-09, 2.92448e-09, -8.011625e-10, 
    6.895107e-11, 8.369945e-10, -8.115713e-10, -6.942749e-10, 5.647678e-09, 
    1.37203e-09, 6.255618e-09, -1.264766e-10, -4.175206e-09, 9.56868e-09, 
    9.56237e-09, -9.757741e-10, -9.063854e-09, 7.715016e-09, 2.116906e-09, 
    -1.191665e-10, 2.819291e-10, 3.34996e-10, -8.469314e-11, -6.405685e-10,
  -8.497523e-10, 2.37327e-09, -5.358061e-10, -4.893081e-10, 5.531433e-10, 
    9.873702e-11, -1.343415e-08, 4.631715e-09, 5.517791e-10, 6.82121e-12, 
    -1.217643e-09, 5.916831e-09, -1.174578e-08, 2.41215e-09, 5.550419e-09, 
    -1.140591e-08, 3.365989e-09, -1.39313e-08, 2.858572e-08, -4.304411e-09, 
    -9.345342e-09, -9.606538e-11, 2.289084e-10, -2.594675e-09, -6.129426e-10, 
    3.355467e-10, 2.595465e-08, 1.627893e-08, 1.577115e-08, -2.385286e-08, 
    1.819961e-08, 1.905482e-08, 2.742405e-08, -1.683702e-10, -9.721418e-09, 
    -1.792478e-08, 5.018023e-10, 1.046722e-09, 1.753449e-08, -3.50548e-09, 
    6.946072e-09, -2.606214e-09, 1.146279e-08, 7.835608e-10, 2.164307e-08, 
    3.47149e-08, 5.670651e-08, 5.956196e-10, -1.390711e-08, -5.432454e-11, 
    -2.082309e-09, -1.105207e-09, 1.368309e-08, -6.054847e-10, -2.220898e-09, 
    3.257981e-10, -1.708804e-08, 4.321469e-08, 1.912323e-08, -1.361092e-08, 
    -8.224788e-09, -5.031552e-09, -1.402896e-10, -1.933165e-09, 
    -5.160189e-09, 5.677691e-09, -2.397377e-08, -1.43545e-08, -1.29819e-09, 
    -7.011806e-09, -1.147043e-09, 2.203217e-08, 2.074785e-11, -3.944365e-10, 
    2.364137e-08, -9.640644e-11, 5.042224e-10, -5.654641e-09, 3.223775e-09, 
    -9.138319e-09, -1.907821e-08, -4.387307e-09, 7.597379e-09, 4.012009e-10, 
    9.154178e-09, -6.93376e-10, -5.24858e-09, -1.180638e-10, 6.389147e-10, 
    -1.226917e-08, 9.633823e-09, 1.373174e-08, -4.364026e-09, -4.146953e-08, 
    -7.85343e-09, -5.736609e-09, -1.720753e-09, -2.534745e-08, 2.737409e-09, 
    -1.110993e-09, -5.486527e-10, 6.873695e-09, -5.888268e-11, -1.016634e-09, 
    -1.073124e-08, 9.723692e-09, 6.317237e-09, -1.08779e-08, -1.886633e-10, 
    6.727817e-09, 3.818343e-09, -2.481386e-09, -1.695071e-09, 1.258775e-08, 
    3.48399e-09, -3.025093e-10, 4.168115e-10, 4.713581e-10, -5.380585e-11, 
    -2.240654e-09,
  -3.515765e-10, 2.842341e-09, -2.684317e-09, -6.042455e-11, 4.393996e-10, 
    -2.996671e-09, -1.674636e-08, 5.536492e-09, 2.630372e-09, 2.439549e-09, 
    -2.605134e-09, 1.659998e-09, -7.118842e-09, 6.259256e-09, 1.562654e-08, 
    -1.754289e-08, 3.315318e-09, -1.897112e-08, 2.894012e-08, -1.502144e-09, 
    -5.387108e-09, -4.532808e-09, -1.561489e-09, -2.092236e-09, 1.728949e-09, 
    2.483318e-09, 4.337255e-08, -1.203944e-10, -1.009084e-08, -2.042179e-08, 
    1.155007e-08, 3.159283e-08, 3.851534e-08, 1.717524e-09, -2.616559e-09, 
    -1.748907e-08, -1.15287e-09, 1.424013e-09, 8.978304e-09, -6.345211e-09, 
    7.876759e-09, -7.357698e-09, 1.425822e-08, 1.364489e-09, 1.805449e-08, 
    1.408654e-08, 7.328393e-08, -3.707896e-10, -1.138508e-08, -1.279545e-10, 
    -2.01134e-09, -9.145992e-09, 1.204004e-08, -1.043566e-09, -6.933861e-09, 
    5.341008e-10, -2.405937e-08, 4.049709e-08, 6.491611e-08, -2.682026e-08, 
    -7.690232e-09, 3.645255e-09, -1.437115e-09, -4.680544e-09, -7.971596e-09, 
    4.947424e-09, -5.285892e-08, -1.36713e-08, -4.824301e-09, -5.661661e-09, 
    -2.610022e-09, 2.133083e-08, -3.04322e-08, 3.616606e-09, 3.199458e-08, 
    1.668923e-10, 5.054162e-10, -8.149215e-09, 5.855492e-09, 1.162164e-08, 
    -3.233163e-08, -5.424498e-09, 4.839109e-09, 5.755396e-10, 2.938179e-09, 
    3.991943e-09, -1.012444e-08, -3.6855e-09, -3.775087e-09, -1.868793e-08, 
    3.681293e-09, 1.221262e-08, -5.999098e-09, -2.190861e-08, -1.478293e-08, 
    -1.910615e-09, -2.194361e-09, -3.68608e-08, 1.635442e-09, -1.645139e-09, 
    -1.219973e-09, 1.314736e-08, 6.993623e-10, -1.071104e-09, -9.884445e-09, 
    5.068841e-09, 1.513285e-09, -1.272832e-08, 5.120171e-09, 5.404672e-09, 
    2.755996e-09, -6.056268e-09, 4.170374e-09, 1.436479e-08, -3.143441e-11, 
    -5.526999e-10, 5.625509e-10, 5.627605e-10, -2.699352e-11, -3.030323e-09,
  1.010164e-09, -1.116405e-10, 3.322782e-09, 6.040921e-09, 1.729347e-09, 
    -2.281638e-09, -9.263829e-09, 2.89981e-09, 9.564019e-09, 1.253738e-09, 
    9.545147e-10, 1.377998e-09, -3.148898e-09, -5.506877e-09, 3.957325e-08, 
    -2.249702e-08, 2.604452e-09, -1.992143e-08, 2.66006e-08, -4.766548e-09, 
    5.435595e-09, -1.418294e-08, -2.71524e-09, 1.877822e-09, 2.549484e-09, 
    3.023843e-09, 5.365558e-08, -2.93187e-09, -9.56548e-08, -1.489008e-08, 
    9.229723e-09, 3.178599e-08, 5.219965e-08, -8.476491e-10, 2.469847e-09, 
    -1.444397e-08, -9.757287e-10, 1.719052e-09, 2.439208e-09, -1.370582e-08, 
    1.252467e-08, -1.269882e-09, 1.68758e-08, 2.233897e-09, 1.875833e-09, 
    -8.55789e-09, 1.041121e-07, -1.005702e-10, -9.208737e-09, -2.224532e-10, 
    -2.396099e-09, -1.582436e-08, 7.749503e-09, -2.881802e-09, -1.550896e-08, 
    6.683933e-10, -4.366308e-08, 3.625482e-08, 1.166669e-07, -1.736167e-08, 
    -4.788035e-09, 8.213419e-09, -1.265562e-09, -9.508529e-09, -1.024285e-08, 
    2.084101e-08, -9.533181e-08, -1.189755e-08, 6.635446e-09, 7.377707e-09, 
    -3.308628e-09, -1.788237e-09, -5.82454e-08, 8.586994e-09, 3.54681e-08, 
    5.289849e-10, 5.837109e-10, -1.138645e-08, 7.410894e-09, 3.982626e-08, 
    -2.971584e-08, 8.966646e-09, 1.838686e-09, 1.729916e-09, -3.381558e-09, 
    7.075812e-09, -6.474352e-09, -6.713378e-09, -1.659494e-09, -3.361404e-08, 
    1.683588e-09, 6.100027e-09, -5.308735e-09, 1.841734e-08, -1.928862e-08, 
    4.912784e-09, -1.852447e-09, -3.001281e-08, -5.880452e-10, -2.75561e-09, 
    -1.890555e-09, 1.132377e-08, 8.864163e-10, -1.20885e-09, 2.369489e-08, 
    -1.013518e-10, -3.992284e-09, 3.28771e-09, 1.312782e-08, 4.512344e-09, 
    1.551939e-09, -5.219704e-09, 4.141441e-09, 1.030122e-08, -7.490144e-09, 
    -9.074256e-10, 9.653007e-10, 6.211796e-10, 1.046274e-11, -5.638299e-09,
  1.110777e-09, -1.814556e-09, 2.947939e-08, 1.728381e-08, 2.736272e-09, 
    -6.693313e-10, 1.017838e-09, -2.09161e-09, 8.133725e-09, 4.437197e-10, 
    2.11179e-09, 9.814585e-10, -5.51438e-10, 4.45084e-11, -1.591167e-08, 
    -2.798559e-08, 1.637454e-09, -2.293501e-08, 2.242713e-08, -4.197261e-09, 
    2.055742e-08, -1.631707e-08, -2.394188e-09, 5.045877e-09, 1.147669e-09, 
    1.995375e-09, 4.125292e-08, 1.213436e-09, -4.336533e-08, -1.341431e-08, 
    2.434234e-08, 4.728668e-08, 6.811092e-08, -8.480242e-09, -1.821263e-09, 
    -1.579502e-08, -1.685083e-09, 2.063778e-09, -2.366676e-08, -1.056247e-08, 
    2.61025e-08, 4.746369e-09, 1.789611e-08, 3.621537e-09, -5.713616e-09, 
    -2.263505e-10, 1.206633e-07, 2.71146e-09, -1.479209e-08, -4.045617e-10, 
    1.081176e-09, -1.072164e-08, 3.72001e-09, -2.072625e-09, -1.070182e-08, 
    5.704521e-10, -3.397349e-08, 3.285565e-08, 1.480454e-07, -2.846303e-08, 
    -9.749158e-09, 6.494474e-09, 4.177366e-09, -1.431416e-08, -9.726454e-09, 
    1.316539e-08, -9.835179e-08, -2.37992e-08, 3.72421e-09, -9.989776e-09, 
    3.710454e-09, -2.635232e-08, -6.930486e-08, 3.867854e-09, 3.966919e-08, 
    8.197958e-10, 1.087386e-09, -1.718044e-08, 5.296453e-09, 3.872958e-08, 
    -3.133817e-08, 3.061238e-08, -1.094065e-09, 2.099569e-09, -1.438252e-09, 
    6.717016e-09, -1.242142e-09, -3.282821e-09, 9.278143e-10, -4.939392e-08, 
    -1.315186e-09, 4.998398e-09, -3.622091e-09, 6.416317e-08, -2.323458e-08, 
    1.911424e-08, 1.931858e-09, -2.37435e-09, -3.8753e-09, -4.416131e-09, 
    -3.277819e-09, 2.925688e-09, 6.256897e-09, -1.236238e-09, 2.438804e-08, 
    -1.138119e-09, -4.179697e-10, 1.124414e-08, 1.414685e-08, 2.814375e-09, 
    -5.362608e-10, -8.784014e-10, 1.990145e-09, 5.22175e-09, -1.929016e-08, 
    -1.513257e-09, 1.653298e-09, 6.137331e-10, 5.286083e-11, -6.449284e-09,
  1.446097e-10, 2.485194e-09, 7.785786e-08, 1.309877e-08, 5.515631e-09, 
    -1.199396e-09, 6.248001e-09, -1.460489e-08, 1.680974e-09, 2.863771e-10, 
    1.611852e-09, 2.413231e-09, 5.346692e-10, 3.412197e-09, -1.330091e-08, 
    -3.165452e-08, -6.588152e-11, -1.32103e-08, 1.706658e-08, 2.716661e-09, 
    2.217826e-08, -2.137085e-09, -7.309836e-09, 9.740575e-09, -3.656169e-10, 
    7.850076e-10, 1.646538e-08, 1.090052e-08, 4.615799e-09, 2.615889e-08, 
    5.662969e-09, 4.976425e-08, 1.012664e-07, -3.223113e-08, -4.969252e-09, 
    -2.108425e-08, -3.397008e-09, 2.27314e-09, -1.74349e-08, -9.991368e-10, 
    4.27096e-08, 5.324637e-09, 1.499933e-08, 4.612897e-09, -1.153467e-08, 
    1.786907e-08, 1.363592e-07, 1.035653e-08, -1.435824e-08, -9.116405e-10, 
    9.413213e-09, -1.785781e-08, -1.780505e-08, -4.435992e-09, -5.688849e-09, 
    2.16005e-10, -2.232616e-08, 3.469735e-08, 1.45459e-07, -4.071026e-08, 
    4.795993e-09, 8.821644e-09, 7.123845e-09, -2.130969e-08, -6.958294e-09, 
    1.105911e-08, -1.083191e-07, -4.07515e-08, 1.593958e-08, -1.561125e-08, 
    1.007186e-08, -4.550691e-08, -6.388279e-08, -4.535309e-09, 5.296137e-08, 
    8.027428e-10, 5.097576e-10, -2.736513e-08, 2.523612e-09, 1.308501e-08, 
    -2.935025e-08, 2.784474e-08, -2.920217e-09, 2.267598e-09, -5.660695e-09, 
    4.722438e-09, 2.187562e-09, 5.254151e-09, 1.064985e-09, -6.101743e-08, 
    -5.888865e-09, 2.397987e-08, -1.502116e-09, 1.484569e-07, -3.164303e-08, 
    4.361326e-08, 1.84825e-08, 1.687067e-08, -6.710593e-09, -5.831862e-09, 
    -2.24918e-09, -5.975025e-10, 9.747978e-09, -7.047234e-10, 2.232548e-08, 
    5.344418e-10, -1.140961e-09, 6.953087e-10, 7.885433e-09, 4.664571e-10, 
    -1.869239e-09, 6.277787e-10, 1.142553e-10, 1.650392e-09, -2.436627e-08, 
    -2.279137e-09, 2.514469e-09, 9.227286e-10, 7.106848e-11, -1.302055e-09,
  3.181589e-08, 5.220102e-09, 9.908644e-08, 5.947811e-09, 7.10935e-09, 
    -6.474068e-09, 6.564676e-09, -1.693667e-08, -4.595393e-09, -1.293131e-09, 
    2.062222e-09, 3.618368e-09, 1.050068e-09, 1.018003e-08, 4.625349e-10, 
    -3.398223e-08, -2.014951e-09, -2.921752e-09, 1.574853e-08, 6.782273e-09, 
    -1.80973e-08, -2.113495e-09, -1.289055e-08, 1.058191e-08, -1.620606e-10, 
    -8.640768e-10, -2.625598e-10, 1.088455e-08, -9.738017e-09, 4.582517e-08, 
    -1.004452e-08, -1.356909e-09, 1.010099e-07, -3.732117e-08, -2.801755e-09, 
    -2.574626e-08, -3.631419e-09, 3.195908e-09, 2.010552e-10, 1.699618e-10, 
    4.557856e-08, 7.98974e-09, 1.622004e-08, 2.152396e-09, 5.236814e-09, 
    1.609425e-08, 1.303791e-07, 2.388967e-08, 9.880717e-09, -1.911282e-09, 
    1.655765e-08, -3.225381e-08, -3.211878e-08, -8.374934e-09, -9.896834e-09, 
    -3.322498e-10, -2.109522e-08, 5.211185e-08, 1.243893e-07, -3.664623e-08, 
    1.770576e-08, 8.519066e-09, 5.767731e-09, -3.147146e-08, -3.34154e-09, 
    2.671271e-08, -4.874738e-08, -5.424494e-08, 2.178621e-08, 4.003726e-08, 
    4.16577e-09, -7.251998e-08, -3.873146e-08, -5.504887e-09, 7.233079e-08, 
    2.531237e-10, -1.331173e-09, -4.184255e-08, 1.625369e-09, 1.592184e-10, 
    -2.905739e-08, 1.922535e-08, -3.213927e-09, 5.286438e-12, -5.275695e-09, 
    -6.567308e-08, 1.278119e-08, 5.355844e-09, 7.863393e-09, -7.89563e-08, 
    -8.565451e-09, 6.089732e-08, -7.534595e-11, 2.367536e-07, -5.091698e-08, 
    5.389307e-08, 4.597452e-08, 1.616166e-08, -8.081031e-09, -6.321022e-09, 
    8.226948e-10, -4.575895e-12, 5.863747e-09, 4.800924e-10, 6.479019e-08, 
    2.623034e-08, -8.228938e-09, -9.724715e-09, 4.460446e-09, -2.28448e-09, 
    -4.35881e-09, 9.659402e-10, -1.31314e-09, -1.966043e-09, -7.858432e-09, 
    -3.188393e-09, 3.255721e-09, 8.578347e-10, 3.313261e-11, 3.676121e-09,
  8.882915e-08, -1.450474e-09, 8.281091e-08, 6.570815e-09, -6.49095e-10, 
    -1.4043e-08, 3.381558e-09, -9.633311e-09, -1.591405e-08, -2.003731e-10, 
    3.308571e-09, 3.545722e-09, 2.640888e-09, 1.174448e-08, 4.047649e-09, 
    -3.652024e-08, -4.842263e-09, 5.642846e-10, 1.899126e-08, -6.473897e-10, 
    -4.534382e-08, -2.155758e-08, 3.088473e-09, 9.749726e-09, -5.147172e-10, 
    -5.983964e-09, 4.769998e-08, 1.790551e-08, -1.259622e-08, 7.40593e-08, 
    -6.831618e-08, -9.896422e-08, 6.016541e-08, -4.259715e-08, -4.242395e-09, 
    -3.6686e-08, -3.204593e-09, 5.136158e-09, 1.557225e-09, 9.174414e-09, 
    3.254305e-08, 9.616144e-09, 1.692075e-08, 4.197176e-11, 2.505942e-09, 
    4.439181e-08, 1.152742e-07, 4.076321e-08, 2.593573e-08, -3.337504e-09, 
    2.514379e-08, -5.661292e-08, -3.36228e-08, -1.040497e-08, -6.317089e-09, 
    -1.003798e-09, -5.860858e-08, 7.71995e-08, 1.103486e-07, -2.866017e-08, 
    7.504411e-09, 4.75967e-09, 4.696801e-09, -4.498228e-08, 1.446358e-09, 
    2.855865e-08, 4.155822e-10, -6.154113e-08, 1.920142e-08, 4.108387e-08, 
    5.084132e-09, -7.094997e-08, -3.320775e-08, 8.787424e-10, 9.890827e-08, 
    -1.217416e-09, -2.072937e-09, -5.9885e-08, 9.463946e-10, -2.035046e-08, 
    -3.331667e-08, 2.102187e-08, -3.170555e-09, -7.581036e-09, 6.823541e-09, 
    -1.036955e-07, -4.668266e-09, 3.821413e-09, 1.425383e-08, -8.614563e-08, 
    -7.096276e-09, 1.219065e-07, 8.526513e-12, 2.825403e-07, -9.875026e-08, 
    5.364207e-08, 2.849405e-08, 9.587723e-09, -7.051369e-09, -8.558425e-09, 
    5.950767e-09, -4.661786e-09, -7.14563e-09, 9.02368e-10, 1.667527e-07, 
    4.600537e-08, -7.707911e-09, -2.053065e-08, -5.884999e-10, -6.444338e-10, 
    -4.803098e-09, 4.229719e-10, -1.096453e-09, -2.023341e-09, 3.668731e-09, 
    -3.856792e-09, 3.240146e-09, 5.55513e-10, -3.698375e-11, 3.558341e-09,
  5.817355e-08, -7.204449e-09, 4.941114e-08, -2.608397e-08, -5.1798e-09, 
    -7.153176e-09, -8.403731e-09, 4.392973e-09, -1.566696e-08, 3.99109e-09, 
    4.397634e-09, 3.023956e-09, 9.929408e-10, -1.626518e-09, 5.084758e-09, 
    -3.909967e-08, -1.675588e-08, -2.520437e-09, 1.647105e-08, -6.88965e-09, 
    -6.252446e-08, -1.538865e-09, -1.927663e-08, -4.234266e-09, 
    -1.463025e-08, -3.232572e-09, 2.452606e-07, 1.193496e-08, 1.02599e-08, 
    7.238441e-08, -2.948548e-08, -1.247436e-07, 3.222567e-09, -1.221156e-08, 
    -2.060222e-08, -5.643949e-08, -3.672199e-10, 7.64139e-09, 3.558648e-08, 
    2.460691e-08, 1.941887e-08, 6.824735e-09, 1.116061e-08, 1.34083e-09, 
    -9.174528e-11, 4.22026e-08, 1.248112e-07, 9.132012e-08, 3.361777e-08, 
    -4.56437e-09, 2.850332e-08, -7.714607e-08, 4.106482e-09, -1.231074e-08, 
    7.837871e-09, -5.085781e-10, -1.083372e-07, 9.507024e-08, 1.05557e-07, 
    -1.295881e-08, 1.8332e-09, 1.482249e-09, 3.480079e-08, -5.521245e-08, 
    7.624704e-09, 2.221259e-08, 3.722243e-08, -7.105496e-08, 1.843728e-08, 
    1.915453e-08, -2.783054e-10, -1.112983e-07, -4.712717e-08, 1.233434e-08, 
    1.280871e-07, -2.726438e-09, -1.673001e-09, -7.336905e-08, -6.487255e-11, 
    3.504852e-09, -3.801597e-08, 2.567074e-08, -2.930165e-09, -9.450105e-09, 
    4.870685e-09, -6.571952e-08, 9.080509e-09, 1.141871e-09, 9.973872e-09, 
    -1.034844e-07, -2.924253e-09, 1.946976e-07, -2.058584e-10, 3.193658e-07, 
    -1.378866e-07, 4.248276e-08, 1.031522e-08, 3.27401e-08, -4.831691e-09, 
    -1.573621e-08, 2.335173e-08, -1.092774e-08, -1.114284e-08, -1.862489e-09, 
    7.304561e-08, 4.213337e-08, -8.278789e-09, -2.816046e-08, -6.749474e-09, 
    4.102958e-10, -3.654577e-09, -8.601546e-10, -3.684818e-09, -8.641337e-10, 
    1.859803e-09, -4.337573e-09, 2.278071e-09, 1.354223e-10, -1.267679e-10, 
    -1.146077e-08,
  -3.439459e-08, -5.094421e-09, 5.517222e-09, -6.453229e-08, -3.377295e-09, 
    9.198175e-09, -1.720468e-08, 1.723788e-08, -1.733156e-09, 5.084871e-09, 
    8.757297e-10, 5.469474e-10, 1.843887e-09, -1.673072e-08, -3.195737e-09, 
    -3.652927e-08, -2.657639e-08, 6.277446e-09, -8.681269e-10, 4.703679e-09, 
    -5.775837e-08, 4.220828e-08, -1.206217e-08, -3.619789e-08, -5.986863e-09, 
    3.729838e-09, 1.571794e-07, -1.353987e-08, 9.847327e-09, 6.840003e-08, 
    2.05489e-08, -6.100231e-08, -1.722685e-08, 2.151978e-08, -3.860237e-08, 
    -6.728067e-08, 3.969285e-09, 8.230657e-09, 4.317337e-08, 4.035858e-08, 
    1.391882e-08, 2.280899e-09, 3.758061e-09, 9.078907e-10, -2.265904e-08, 
    1.199999e-08, 1.240143e-07, 1.559652e-07, 3.577379e-08, -5.284939e-09, 
    3.335943e-08, -5.449886e-08, 6.307508e-08, -1.122269e-08, 2.013479e-08, 
    -1.20906e-10, -1.537694e-07, 1.030864e-07, 8.17619e-08, 8.149485e-09, 
    1.431658e-09, 3.013838e-10, 5.441154e-08, -4.635149e-08, -1.483979e-08, 
    1.907392e-08, 5.623679e-08, -6.593768e-08, 1.274589e-08, 3.837249e-08, 
    2.021682e-08, -1.422999e-07, -5.4515e-08, 9.952714e-09, 1.407611e-07, 
    -1.735089e-09, 1.572033e-09, -7.819202e-08, -5.419224e-10, -6.808807e-08, 
    -4.174228e-08, 2.916948e-08, -3.904972e-09, -3.97813e-09, 5.118181e-10, 
    -5.69953e-08, 2.916136e-08, -4.053504e-09, 9.854618e-09, -1.161713e-07, 
    -2.017146e-09, 2.650305e-07, -4.228298e-10, 3.797223e-07, -7.827498e-08, 
    3.045295e-08, -2.95779e-08, 6.25563e-08, -6.630557e-09, -2.492375e-08, 
    -2.199499e-09, -4.610357e-09, -1.335558e-08, -4.036281e-09, 
    -3.586217e-08, 2.810805e-08, -8.276288e-09, -2.89624e-08, -7.330755e-09, 
    2.626166e-10, -1.568878e-11, 6.65068e-11, -4.859203e-09, -8.049028e-10, 
    -1.828312e-09, -4.540743e-09, 8.942607e-10, -4.016698e-10, -2.077698e-10, 
    -1.539001e-08,
  -7.349263e-08, -1.176431e-09, -2.299771e-09, -4.02058e-08, 1.112812e-08, 
    1.597346e-08, -1.266835e-08, 2.062166e-09, 2.471256e-08, 2.003617e-09, 
    -1.538183e-10, -4.069989e-11, 1.546869e-08, -2.383786e-08, -1.577098e-08, 
    -3.85855e-08, -4.665723e-08, 2.03836e-08, -4.847216e-08, 2.080719e-08, 
    -4.662263e-08, 7.044252e-08, 3.676496e-08, -1.030912e-09, 1.024966e-08, 
    3.95903e-09, 2.985712e-08, -1.161857e-08, 1.049216e-08, 7.938786e-08, 
    3.470586e-08, -2.114143e-08, -1.434296e-08, -2.661295e-09, -5.176958e-08, 
    -8.71853e-08, 8.819654e-09, 9.427069e-09, 3.506386e-08, 5.096994e-08, 
    -3.371838e-08, 3.394007e-09, 2.439151e-10, -1.210626e-09, -3.180094e-08, 
    -1.949979e-08, 7.767676e-08, 2.008135e-07, 3.608775e-08, -5.199631e-09, 
    3.806996e-08, -4.196204e-08, 1.700688e-07, -1.265321e-08, 3.491184e-08, 
    -6.838832e-10, -1.599948e-07, 1.028486e-07, 6.14907e-08, 1.299455e-08, 
    -3.001333e-11, 2.098659e-10, -9.605969e-09, -2.464972e-08, -9.815474e-08, 
    1.855688e-08, 2.904324e-08, -8.009647e-08, 3.669811e-09, 5.414188e-08, 
    4.693555e-07, -1.363082e-07, -7.311576e-08, 4.107278e-09, 1.371515e-07, 
    -2.881961e-10, 3.345733e-09, -7.038665e-08, -5.078704e-10, -1.22907e-07, 
    -4.818367e-08, 4.27866e-08, -1.416879e-08, -1.811031e-09, -5.126594e-09, 
    -3.338232e-08, -1.021988e-08, -5.526886e-09, 1.400273e-08, -1.226571e-07, 
    9.601422e-09, 2.999317e-07, -1.837236e-09, 4.172621e-07, -4.98834e-08, 
    1.934818e-08, -3.584707e-08, 3.318564e-08, -1.838748e-08, -3.403332e-08, 
    -4.009905e-08, 6.529262e-09, -1.132477e-08, -1.788516e-08, -3.324919e-08, 
    1.576382e-08, -1.965452e-08, -1.759815e-08, -2.231786e-09, -1.504532e-09, 
    4.34045e-09, -2.482921e-10, -4.095114e-09, -3.205287e-09, -1.147669e-09, 
    -4.381036e-09, -7.70342e-10, -6.614194e-10, -2.983924e-10, -3.291689e-09,
  -4.813688e-08, 1.064279e-09, 1.644713e-08, 1.110203e-08, 1.273662e-08, 
    9.714483e-09, 9.96863e-10, -6.9154e-09, 1.283621e-08, 4.826006e-11, 
    -1.313936e-09, 8.845404e-10, 3.018243e-08, -3.014742e-08, -6.893686e-09, 
    -3.867283e-08, -5.263497e-08, 5.170097e-08, -1.859803e-07, 2.994767e-08, 
    -3.797567e-08, 4.337079e-08, 6.424585e-08, 1.776783e-08, 8.717336e-09, 
    7.649419e-10, -6.147786e-09, -5.809227e-09, 7.86639e-09, 9.00821e-08, 
    9.535881e-09, -2.54164e-09, -6.212815e-09, 1.3906e-08, -6.713111e-08, 
    -1.182296e-07, 9.572659e-10, 1.249603e-08, 1.894722e-08, 3.817847e-08, 
    -1.582059e-07, 7.244523e-09, -5.024674e-10, -4.368907e-09, -3.31583e-08, 
    -4.794987e-08, 1.101115e-07, 2.332941e-07, 3.938013e-08, -4.605425e-09, 
    4.162553e-08, -4.03341e-08, 2.454251e-07, -1.62125e-08, 5.614859e-08, 
    -2.496279e-09, -1.420531e-07, 8.705454e-08, 7.039169e-08, 7.462802e-09, 
    2.032152e-10, -3.282372e-08, 4.60858e-09, -1.147445e-08, -1.528678e-07, 
    3.158692e-08, 3.879762e-08, -9.469107e-08, -5.613344e-09, 5.796272e-08, 
    2.833534e-07, -7.630143e-08, -1.00189e-07, 7.159031e-09, 1.439813e-07, 
    -5.573668e-09, 5.457409e-09, -6.081194e-08, -1.962746e-10, -8.191597e-08, 
    -5.637992e-08, 7.15769e-08, -4.041721e-08, -2.142428e-10, -2.247077e-09, 
    -4.192714e-09, -8.817682e-08, -4.544916e-09, 2.637329e-08, -9.795406e-08, 
    4.916654e-08, 2.642734e-07, -3.992824e-09, 4.125282e-07, -4.735699e-08, 
    7.233052e-09, -5.197161e-08, -1.936422e-08, -2.009682e-08, -4.290092e-08, 
    -1.264808e-07, 4.970182e-09, -2.566807e-09, -2.651743e-08, -4.42447e-08, 
    4.112434e-08, -1.622999e-08, -7.262486e-09, -6.974119e-10, 3.933621e-09, 
    4.375181e-09, -2.623949e-09, -7.564665e-09, -9.597841e-09, 1.032845e-10, 
    -3.782407e-09, -7.701573e-10, -6.646026e-10, -4.246914e-10, -4.535383e-08,
  -3.491488e-08, 2.353715e-09, 2.740438e-08, 2.399764e-08, 8.69835e-09, 
    1.594054e-08, 2.560176e-08, -2.696419e-08, -6.702351e-09, -4.718515e-09, 
    -2.343143e-09, -1.109299e-09, 2.121834e-08, -3.350863e-09, -1.381471e-08, 
    -3.616634e-08, -4.78111e-08, 7.864071e-08, -3.023912e-07, 2.603036e-08, 
    -2.542328e-08, 4.582256e-08, 4.400255e-08, 4.881315e-09, -9.066525e-11, 
    -2.781405e-09, -1.35588e-08, -4.660194e-09, 2.182713e-08, 8.632691e-08, 
    8.953691e-09, 4.175774e-09, -1.627939e-09, 1.033807e-07, -9.173328e-08, 
    -1.528663e-07, -1.799037e-09, 1.844928e-08, 1.394352e-08, 1.151389e-08, 
    -2.316319e-07, 6.451558e-09, -4.046882e-09, -5.368555e-09, -7.415736e-09, 
    -6.501529e-08, 1.52845e-07, 2.13755e-07, 3.389197e-08, -4.093096e-09, 
    4.469914e-08, -3.261113e-08, 2.837771e-07, -1.603938e-08, 8.061075e-08, 
    -6.994014e-10, -1.332357e-07, 6.142626e-08, 9.362966e-08, -1.686263e-08, 
    1.918863e-09, -9.953675e-08, 1.362451e-08, -2.126566e-08, -8.209601e-08, 
    7.678642e-08, -1.183486e-08, -9.183765e-08, -1.331449e-08, 3.931729e-08, 
    -2.087763e-07, -1.538723e-08, -7.881869e-08, 4.556057e-09, 1.814986e-07, 
    -1.816414e-08, 1.027573e-08, -3.336788e-08, 5.386755e-09, -5.514534e-08, 
    -5.233494e-08, 1.151235e-07, -5.551357e-08, -1.536534e-09, -2.317677e-09, 
    -7.796814e-09, -2.042579e-07, 1.103803e-08, 4.869478e-08, -1.531289e-07, 
    7.092609e-08, 1.801294e-07, -4.712547e-09, 3.921678e-07, -9.393926e-08, 
    -1.097226e-08, -3.245314e-08, 7.259757e-09, -3.234157e-08, -5.07827e-08, 
    -1.415853e-07, -1.823065e-08, -4.687593e-10, -2.774198e-08, 
    -7.587397e-08, 7.833404e-08, 7.941537e-09, -1.037125e-08, 4.732613e-09, 
    3.301426e-08, 9.112e-11, -4.560377e-09, -1.206234e-08, -1.773248e-08, 
    -6.543871e-09, -3.035211e-09, 1.534943e-09, -7.51065e-10, -5.518856e-10, 
    -6.78985e-08,
  -2.48192e-08, 5.911943e-09, 9.69851e-09, 1.837941e-08, 1.467231e-08, 
    1.858928e-08, 4.297362e-08, -2.41339e-08, -2.641286e-08, -1.434955e-08, 
    3.275773e-09, -1.66051e-09, -2.340141e-08, 7.826088e-09, -6.720143e-09, 
    -3.148096e-08, -5.201991e-08, 6.960147e-08, -2.549475e-07, -1.885542e-08, 
    8.474785e-09, 1.769967e-07, 2.057266e-08, -1.893909e-09, -2.285128e-08, 
    -1.279132e-07, -3.650598e-09, -1.298008e-08, 2.89109e-08, 9.168389e-08, 
    1.674277e-08, 1.899718e-08, -1.320927e-09, 1.197874e-07, -1.392939e-07, 
    -1.222347e-07, -1.06797e-08, 2.556315e-08, 3.053424e-08, 7.275851e-10, 
    -2.379113e-07, 3.444825e-09, -1.021715e-08, -4.991723e-09, -1.854585e-08, 
    -6.720688e-08, 1.319942e-07, 1.259613e-07, -1.01357e-08, -6.863445e-09, 
    4.715524e-08, -3.99873e-08, 2.302032e-07, -1.68081e-08, 1.125652e-07, 
    -5.641198e-09, -1.47396e-07, -3.835726e-08, 1.086177e-07, -1.77473e-08, 
    2.51805e-09, -9.301209e-08, -7.726908e-08, -3.225057e-08, -4.931515e-08, 
    7.205631e-08, 7.752533e-09, -1.03413e-07, -2.167837e-08, 3.248726e-08, 
    -2.873113e-07, 5.846186e-08, -9.42789e-08, -1.316039e-09, 1.81514e-07, 
    -2.910554e-08, 1.264171e-08, -2.255518e-09, 1.591835e-08, -7.355766e-08, 
    -3.938459e-08, 1.352734e-07, -3.535035e-08, -8.060579e-08, -6.815822e-08, 
    -2.988895e-08, -3.370656e-08, 3.494165e-08, 7.073768e-08, -1.71546e-08, 
    3.082187e-08, 9.995367e-08, -5.43227e-09, 3.53634e-07, -9.392033e-08, 
    -8.494624e-08, 2.125805e-08, 1.370302e-08, -5.127538e-08, -5.550066e-08, 
    -2.033172e-07, -4.826066e-08, -5.180567e-11, -2.066498e-08, 
    -7.630149e-08, 5.204936e-08, -3.763716e-09, -1.264743e-08, 1.779767e-08, 
    6.118682e-08, -2.043407e-09, -2.850243e-09, -1.259582e-08, -2.731531e-08, 
    -8.826078e-09, -2.694185e-09, 7.778937e-09, -7.142837e-10, -6.606697e-10, 
    -5.273466e-08,
  -1.598676e-08, 1.415549e-08, -7.582344e-09, 9.840164e-09, 2.228705e-08, 
    2.591617e-08, 5.689981e-08, -1.828619e-08, -1.691672e-08, -3.593789e-08, 
    -1.927992e-08, -2.517697e-08, -3.593345e-08, -4.940739e-08, 
    -1.304306e-08, -3.266708e-08, -5.300427e-08, 4.189519e-08, -1.555586e-07, 
    -1.093871e-07, 7.60474e-08, 5.583559e-08, 1.277033e-08, -1.486796e-09, 
    -6.544349e-08, -1.48197e-07, 2.462571e-09, -1.448279e-08, 3.103514e-08, 
    1.50001e-07, 2.178342e-08, 9.702489e-09, -5.635798e-09, 1.481183e-07, 
    -1.52916e-07, -5.187485e-08, -1.953501e-08, 2.941846e-08, 3.82405e-08, 
    6.589644e-10, -1.089705e-07, 2.651518e-09, 8.960228e-10, 2.793252e-09, 
    -2.52179e-08, -8.08468e-08, 1.252868e-07, 4.981405e-08, -4.048761e-08, 
    -1.106535e-08, 4.800214e-08, -3.180105e-08, 1.429436e-07, -1.22549e-08, 
    1.271193e-07, -5.192362e-09, -1.617747e-07, 6.01339e-08, 1.096957e-07, 
    -2.206636e-08, 4.964704e-10, -5.264349e-08, -3.418438e-08, -2.841996e-08, 
    -3.445077e-08, 6.222717e-08, 1.205865e-08, -8.932989e-08, -3.174785e-08, 
    2.679462e-08, -1.729037e-07, 7.120047e-08, -1.03261e-07, -5.943321e-09, 
    1.564997e-07, -3.382775e-08, 6.89522e-09, 4.188851e-08, 3.06732e-08, 
    2.598605e-07, -2.768979e-08, 1.2474e-07, 6.405457e-09, -1.319763e-07, 
    -9.925247e-08, -9.908035e-08, 2.694026e-08, 5.793424e-08, 7.581085e-08, 
    -1.17285e-09, -7.584049e-10, 2.888073e-08, -5.256709e-09, 2.976595e-07, 
    -1.066857e-07, 5.20103e-08, 2.786792e-08, 8.412826e-12, -6.466757e-08, 
    -5.197694e-08, -1.131531e-07, -5.044281e-08, -9.174883e-10, 
    -1.389402e-08, -2.170918e-08, -5.004154e-09, -3.38166e-08, -2.180741e-09, 
    2.02017e-08, 5.826291e-08, -9.408154e-09, -1.791022e-09, -8.304937e-09, 
    -3.494324e-08, -4.826347e-09, -1.587307e-09, 1.615835e-08, -5.242065e-10, 
    -7.953957e-10, -4.284163e-08,
  -1.481482e-08, 3.086501e-08, -1.152006e-08, 4.564356e-09, 4.702741e-08, 
    3.932831e-08, 5.88098e-08, -3.102002e-09, 9.040889e-09, -3.557096e-08, 
    -2.657401e-08, -8.780586e-08, -7.089e-09, -6.475585e-08, 6.641869e-09, 
    -5.735507e-08, -4.490436e-08, 2.380909e-08, -7.90378e-08, -4.530608e-08, 
    -5.565204e-08, -2.743315e-08, 1.138837e-07, 3.3628e-09, -8.07525e-08, 
    -1.132418e-07, 1.375855e-08, -1.043833e-08, 2.850282e-08, 2.246862e-07, 
    1.849054e-08, -8.45165e-09, 1.302107e-08, 5.01864e-07, -1.346113e-07, 
    -2.604264e-08, -2.60102e-08, 3.138607e-08, 5.411238e-08, 1.66831e-08, 
    -2.500074e-08, -9.201671e-08, -1.720227e-08, 1.74757e-08, 4.864489e-09, 
    -8.43965e-08, 7.85173e-08, 4.223503e-08, -5.056376e-08, -1.129431e-08, 
    4.72742e-08, -5.928445e-08, 7.858402e-08, -1.539071e-08, 1.236794e-07, 
    -4.596075e-09, -1.770066e-07, 1.555126e-07, 1.095623e-07, -4.898476e-08, 
    -1.431374e-09, -4.988459e-08, 1.300854e-07, 3.984802e-09, -1.59289e-08, 
    3.703786e-08, 1.625193e-08, -7.471527e-08, -3.31267e-08, 1.435689e-08, 
    -5.742714e-08, 2.902993e-10, -4.854479e-08, -4.437254e-09, 1.184632e-07, 
    -3.118583e-08, -1.913406e-09, 6.894351e-08, 2.203674e-08, -1.647227e-07, 
    -2.087273e-08, 8.415267e-08, 3.408405e-08, -1.047781e-07, -5.591534e-08, 
    -5.728003e-08, -5.154101e-08, 6.250008e-08, 7.847824e-08, -6.683575e-08, 
    2.043936e-08, 5.059122e-09, -5.235023e-09, 1.979336e-07, -9.005754e-08, 
    1.027652e-07, 1.252514e-08, -2.248561e-08, -7.175385e-08, -4.900099e-08, 
    -8.228636e-08, -4.139853e-08, -2.666781e-09, -8.069208e-09, 
    -2.494346e-09, -3.254553e-08, -6.01687e-08, 8.135032e-09, 1.053382e-08, 
    3.573501e-08, -4.558018e-08, -1.629985e-09, -5.782283e-09, -3.971826e-08, 
    -1.092587e-09, -1.033561e-09, 2.110353e-08, -8.176499e-10, -9.58174e-10, 
    -8.80645e-08,
  -9.302369e-09, 5.10567e-08, 1.216341e-08, 1.787214e-09, 5.33858e-08, 
    5.208466e-08, 6.66717e-08, 1.120253e-08, 3.566623e-08, -1.531538e-08, 
    -5.304054e-08, -5.929832e-08, 2.801784e-08, -3.584489e-09, 1.834456e-08, 
    -7.162723e-08, -3.810628e-08, 1.375116e-08, -6.097795e-08, 2.069538e-08, 
    2.458165e-08, -4.116265e-08, -7.381328e-08, -4.793577e-08, -6.323484e-08, 
    -7.832017e-08, 3.534086e-08, -1.771338e-08, 1.782024e-08, 2.329107e-07, 
    2.121141e-08, -1.799111e-08, -8.806467e-09, 5.844658e-07, -1.178096e-07, 
    3.623043e-07, -2.708077e-08, 3.17345e-08, 6.124577e-08, 1.649705e-08, 
    2.49741e-08, -2.615674e-07, -9.560779e-08, 3.839169e-08, -9.187431e-09, 
    -7.853754e-08, 1.040065e-07, 8.319677e-08, -4.597413e-08, -7.690744e-09, 
    4.465099e-08, -1.642363e-07, 7.222112e-08, -1.602444e-08, 1.073345e-07, 
    -3.556522e-09, -1.758737e-07, 1.620389e-07, 1.550131e-07, -9.470681e-08, 
    -1.39778e-10, -1.775419e-08, 2.896225e-07, -1.743103e-08, 3.583708e-08, 
    3.366455e-08, 1.985683e-08, -5.32861e-08, -4.398538e-08, -1.828124e-08, 
    4.680129e-08, -9.210731e-08, -2.424377e-08, 7.116284e-09, 8.197192e-08, 
    -2.124438e-08, -1.261495e-08, 7.95537e-08, 2.867258e-08, 2.313101e-08, 
    -6.643972e-09, 5.486651e-08, 5.632762e-08, -7.786963e-08, 1.573664e-07, 
    -4.188809e-08, -1.192321e-07, 3.309191e-08, 5.014591e-08, -1.220627e-07, 
    5.651219e-08, 1.520004e-09, -6.262269e-09, 1.215746e-07, -5.013004e-08, 
    7.605773e-08, -3.876336e-08, -1.231399e-09, -7.881346e-08, -6.696081e-08, 
    -1.350222e-07, -2.650244e-08, -5.336169e-09, -7.70882e-10, 2.459558e-09, 
    -1.558834e-08, -4.335988e-08, 4.044801e-08, -1.014888e-08, 1.287532e-08, 
    -6.699298e-08, -5.592085e-09, -4.680544e-09, -3.894826e-08, -1.93308e-08, 
    1.594708e-09, 1.95855e-08, -1.738396e-09, -1.228216e-09, -1.334672e-07,
  2.647027e-09, 4.90939e-08, 6.334841e-08, 2.606214e-09, 9.675716e-09, 
    3.484678e-08, 7.057855e-08, 1.630116e-08, 5.352985e-08, 1.050154e-08, 
    -5.049577e-08, -2.070061e-08, 2.331939e-08, 4.615327e-08, -1.01416e-08, 
    -6.943534e-08, -2.207508e-08, 4.33505e-08, -4.885496e-08, 1.997017e-08, 
    5.633484e-08, -5.06098e-08, -1.007025e-07, -6.603108e-08, 7.022078e-08, 
    -3.123995e-08, 2.064093e-08, -3.118492e-08, 1.063887e-08, 2.3335e-07, 
    3.371082e-08, -8.959717e-09, -1.641985e-08, 4.213651e-07, -1.364381e-07, 
    4.238103e-07, -2.561676e-08, 2.992611e-08, 4.922214e-08, 3.429841e-08, 
    3.711279e-08, -1.079493e-07, -1.461535e-07, 5.580424e-08, -3.577151e-08, 
    -5.60097e-08, 1.2262e-07, 1.35769e-07, -3.687083e-08, -4.477876e-09, 
    4.075497e-08, -2.427343e-07, 1.212843e-07, -1.814452e-08, 8.259171e-08, 
    -2.053014e-09, -2.017271e-07, 1.261842e-07, 1.261629e-07, -7.303062e-08, 
    -1.752085e-09, 1.1294e-07, -5.462238e-08, -6.777519e-08, 2.461471e-08, 
    3.623626e-08, 1.322843e-08, -5.412136e-08, -3.283657e-08, -4.369832e-08, 
    5.888234e-08, -9.9435e-08, -3.744452e-08, 1.461336e-08, 4.694248e-08, 
    -1.266829e-08, -1.616307e-08, 8.152628e-08, 7.870963e-09, 5.591465e-08, 
    5.163002e-08, 3.717731e-08, 4.123063e-08, -6.329816e-08, 4.671909e-08, 
    -6.350939e-08, -1.788931e-07, 1.322218e-08, 1.686286e-08, -2.181162e-07, 
    5.896783e-08, 1.477237e-08, -8.547147e-09, 8.185492e-08, 1.512564e-08, 
    8.471236e-09, -8.598712e-08, 1.280417e-07, -9.376896e-08, -8.488538e-08, 
    -1.750497e-07, -4.544304e-09, -6.780887e-09, 2.613127e-09, 1.651171e-08, 
    -2.347696e-08, -3.001617e-09, 3.505846e-08, -3.398037e-08, -2.046193e-09, 
    -4.805833e-08, -3.973975e-08, -8.476093e-09, -3.564782e-08, 
    -1.220923e-08, 3.42003e-09, 1.531299e-08, -2.58434e-09, -1.416971e-09, 
    -9.167678e-08,
  -5.62909e-09, 1.808735e-08, 7.943208e-08, 4.951971e-09, -4.053459e-08, 
    -1.033413e-08, 6.723803e-08, 1.904937e-08, 6.166533e-08, 1.422229e-07, 
    -1.593321e-08, 1.757644e-08, 1.918845e-07, 6.231448e-08, -3.738887e-08, 
    -4.963361e-08, -5.181437e-09, 1.179285e-08, -4.574815e-09, -4.67021e-08, 
    3.938226e-08, -2.170805e-08, 5.826564e-08, -3.937589e-08, -1.443266e-07, 
    6.069422e-08, 7.982862e-09, -2.094407e-08, 8.454663e-09, 2.61748e-07, 
    3.20872e-08, 4.59363e-09, -2.632714e-08, 2.803861e-07, -1.273033e-07, 
    3.839357e-07, -2.275074e-08, 2.648886e-08, 9.551286e-09, 4.437513e-08, 
    2.829606e-08, -7.792664e-08, -1.155809e-07, 6.407848e-08, 5.51322e-08, 
    -3.459741e-08, 1.294034e-07, 1.714201e-07, -3.029313e-08, -8.686669e-10, 
    3.559191e-08, -2.291979e-07, 1.82842e-07, -2.066922e-08, 5.084025e-08, 
    -1.107651e-09, -1.612336e-07, 1.146597e-07, 1.514305e-07, -2.60076e-08, 
    -3.303967e-08, 2.268075e-08, -4.559365e-08, -1.701696e-08, 1.013077e-08, 
    3.051105e-08, 2.905381e-09, -5.23894e-08, -3.240211e-08, -3.667083e-08, 
    4.240451e-08, -6.571281e-08, -4.137632e-08, 9.307541e-09, 3.359864e-08, 
    -2.161778e-08, 1.279773e-09, 6.471168e-08, 5.374437e-09, -6.538198e-08, 
    6.445555e-08, 4.793759e-08, 1.981493e-08, -6.740515e-08, -1.282679e-07, 
    -9.498558e-08, -2.004685e-07, -1.470426e-09, -7.974702e-09, 
    -2.439845e-07, 1.37368e-07, 2.785809e-08, -8.119969e-09, 6.369237e-08, 
    3.43648e-08, 6.687375e-08, -1.271437e-07, 4.975914e-08, -1.038791e-07, 
    -6.785026e-08, -1.010937e-07, -1.383314e-07, -9.559216e-09, 3.547584e-09, 
    -2.14709e-09, -5.197398e-08, 3.972445e-08, 5.741185e-09, -4.61132e-08, 
    -1.160379e-08, -3.497939e-08, -6.547589e-08, -2.089496e-08, 
    -3.990749e-08, 5.645006e-09, 3.541595e-09, 1.280443e-08, -2.447038e-09, 
    -1.463107e-09, 1.937224e-09,
  -1.766733e-08, -4.416449e-09, 2.327982e-08, -9.231655e-09, -5.159819e-08, 
    -5.874716e-08, 1.079246e-08, -3.08068e-08, 6.03514e-08, -6.832914e-08, 
    -3.881672e-08, 7.16355e-08, 1.028383e-07, 3.228655e-08, -5.859175e-08, 
    -2.6119e-08, 1.760242e-08, -1.250271e-08, -6.89048e-08, -5.82167e-08, 
    3.255633e-08, 1.646873e-08, 8.428782e-08, -7.166989e-09, -1.021527e-07, 
    2.310441e-07, 3.345161e-08, -1.133043e-08, 3.775824e-09, 1.625825e-07, 
    3.101178e-08, 8.767927e-09, -4.08499e-08, 1.775044e-08, -1.165435e-07, 
    3.14504e-07, -1.860662e-08, 2.392153e-08, -1.15989e-09, 7.01845e-08, 
    -9.787539e-09, -7.342629e-08, -2.132762e-08, 3.54552e-08, -5.025896e-08, 
    -2.841006e-08, 9.088586e-08, 1.912693e-07, 6.932204e-09, 2.344223e-09, 
    2.970772e-08, -1.512361e-07, 2.358377e-07, -1.473937e-08, 1.550814e-08, 
    -2.340926e-09, -1.378059e-07, 1.370502e-07, 8.47671e-08, 1.061454e-08, 
    -3.361939e-07, -4.400539e-08, -1.748134e-08, -1.013349e-08, 
    -4.562984e-08, 3.31425e-08, 2.479226e-09, -3.139218e-08, -2.763881e-08, 
    -1.705047e-08, 6.061515e-08, -3.218537e-08, 7.091614e-09, 2.244741e-08, 
    3.175711e-08, -4.323607e-08, 1.490446e-08, 4.306256e-08, 8.378631e-10, 
    -1.03196e-07, 3.87783e-08, 5.576256e-08, 2.138506e-08, -9.666525e-08, 
    -1.144336e-07, 5.172416e-08, -1.189836e-07, -8.11059e-09, -1.427906e-08, 
    -2.433809e-07, -9.500235e-08, 2.503315e-08, -1.398834e-08, 8.467851e-08, 
    1.309577e-07, 1.903e-07, -1.438427e-07, -5.39444e-11, -1.109457e-07, 
    -9.538861e-08, -2.04181e-08, -5.699388e-08, -1.314811e-08, 4.535075e-09, 
    -1.179063e-08, -5.899375e-08, 3.89262e-08, -1.645316e-08, -4.563498e-08, 
    -1.281825e-08, -3.156771e-08, -5.053136e-08, -5.819862e-08, 
    -3.343706e-08, 4.032756e-09, 2.247236e-09, 1.181371e-08, -2.786514e-09, 
    -1.416666e-09, 4.909379e-08,
  -9.501446e-08, 9.327209e-09, -2.704746e-08, -2.879096e-08, -6.81955e-08, 
    -1.689375e-07, -6.067091e-08, -6.765288e-08, 4.836068e-08, -3.078071e-09, 
    -3.276227e-08, -9.446444e-08, 1.711935e-07, -4.109427e-08, 1.974769e-07, 
    -1.61472e-08, 2.402859e-08, -2.126342e-09, -1.766667e-07, -4.622257e-08, 
    -1.666103e-08, 1.883609e-08, -1.363985e-07, 7.598896e-08, 3.51431e-08, 
    -2.505249e-08, 7.702874e-08, -3.838295e-09, -1.299384e-08, 1.090708e-07, 
    3.286755e-08, -2.44961e-09, -4.286073e-08, -1.789965e-08, -7.027847e-08, 
    2.612409e-07, -2.272428e-08, 2.384391e-08, 1.657099e-08, 7.843472e-08, 
    -7.385413e-08, 1.115459e-07, 5.968172e-08, 4.105888e-08, -4.933474e-08, 
    -3.063735e-08, 8.169087e-08, 1.90253e-07, 4.309575e-08, 3.184198e-09, 
    2.490044e-08, -7.253061e-08, 2.613595e-07, 2.676347e-09, -4.255472e-09, 
    -2.368779e-09, -1.141135e-07, 3.700423e-08, 5.97642e-08, -6.101018e-08, 
    -3.217061e-07, -6.508162e-08, -5.692323e-08, 5.392465e-09, -4.724018e-08, 
    7.10736e-08, -7.18353e-09, -3.448793e-08, -2.799209e-08, -2.495528e-08, 
    3.142213e-08, -8.336201e-09, 1.953936e-08, 2.345967e-07, 9.794974e-09, 
    -2.48383e-08, 4.141228e-09, 5.401461e-08, 1.619535e-08, -1.42029e-08, 
    2.80283e-08, 4.512775e-08, 2.280103e-08, -1.13947e-07, -1.30533e-08, 
    3.933474e-08, -7.044878e-08, -1.511205e-08, -3.525761e-08, -2.290525e-07, 
    -3.456296e-08, 2.080142e-08, -1.242054e-08, 6.740942e-08, 3.293621e-09, 
    9.186234e-08, -1.575582e-07, -1.033072e-08, -8.836719e-08, -8.654663e-08, 
    -1.934632e-08, 7.895038e-08, -1.559109e-08, 5.872955e-09, 1.747787e-08, 
    -6.646508e-08, 1.03214e-08, -3.346861e-08, -3.68849e-08, -1.070214e-08, 
    -2.929403e-08, -2.8714e-08, -5.431264e-08, -1.04767e-08, 3.927425e-09, 
    6.298137e-10, 1.084774e-08, -2.925532e-09, -1.320899e-09, 7.3058e-08,
  -2.76125e-07, 6.130847e-08, 5.093966e-09, -2.5752e-08, -1.964928e-07, 
    -2.453902e-07, -6.784205e-08, -5.079357e-08, 4.389142e-08, -1.820126e-10, 
    -3.625712e-08, -9.206644e-08, -2.164222e-08, 2.218792e-08, -3.023081e-08, 
    -2.545235e-10, 2.054207e-08, 3.576588e-09, -1.556424e-07, -9.306291e-09, 
    7.689891e-09, 2.430113e-08, -2.613298e-07, 1.145747e-08, 3.291018e-08, 
    -9.204075e-08, 9.00335e-08, 9.896439e-10, -1.211367e-08, 1.455206e-07, 
    3.298771e-08, -7.96706e-09, -3.424782e-08, -1.550198e-07, -4.282015e-09, 
    2.249097e-07, -4.1819e-08, 2.599441e-08, 1.292358e-08, 7.590204e-08, 
    -1.186462e-07, 6.409834e-08, 2.912657e-09, 2.191878e-08, -1.065094e-07, 
    -3.01842e-08, 9.841028e-08, 1.648905e-07, 1.560306e-09, 2.455465e-09, 
    2.165558e-08, -7.137908e-08, 2.491383e-07, 1.71425e-08, -2.116789e-08, 
    -2.642992e-09, -1.170725e-07, 3.97101e-09, -6.29416e-08, -8.937508e-08, 
    2.820218e-08, -3.312164e-08, -2.377521e-08, 2.917751e-08, -4.092824e-08, 
    2.864965e-08, -1.881631e-09, -1.373348e-08, -2.758213e-08, 1.707838e-08, 
    7.457515e-09, 2.327283e-09, 1.953254e-09, -1.174919e-08, 7.672316e-09, 
    -8.636903e-09, 7.128705e-09, 5.238621e-08, 4.139145e-08, 5.703657e-08, 
    1.196145e-08, 3.335921e-08, 2.7076e-08, -8.48371e-08, 1.859269e-08, 
    3.203028e-07, -2.859645e-08, -3.06203e-08, -5.520004e-08, -2.082951e-07, 
    -4.509218e-08, 2.511076e-08, -9.300152e-09, 3.877878e-08, -4.50749e-08, 
    4.334502e-08, -2.284332e-07, -2.13073e-08, -7.548658e-08, -4.050865e-08, 
    -6.204834e-08, 6.224944e-08, -1.286992e-07, 6.664251e-09, 1.299406e-08, 
    -6.406515e-08, -8.20171e-09, -4.979177e-08, -3.158254e-08, -7.823814e-09, 
    -2.832724e-08, -1.879687e-08, -1.39961e-08, -2.513275e-09, 3.622404e-09, 
    -7.063136e-10, 1.009047e-08, -2.524445e-09, -1.228159e-09, 1.231035e-08,
  -3.93689e-07, 2.177134e-07, 5.437093e-07, -2.443278e-08, -2.199085e-07, 
    -1.054956e-07, -3.280195e-08, -4.590606e-08, 7.913434e-08, -2.305319e-08, 
    -1.337764e-08, 3.579544e-09, -1.779831e-07, -3.803052e-09, 7.327492e-08, 
    3.337765e-08, -7.990514e-09, 9.498024e-09, -1.026701e-07, 1.082616e-07, 
    1.665626e-08, 1.396677e-08, -1.081854e-07, 1.069589e-08, 4.11859e-08, 
    -6.204652e-08, 9.853534e-08, 6.765276e-09, 2.067077e-08, 1.540177e-07, 
    3.771174e-08, -2.316938e-10, -2.23738e-08, -3.10602e-07, 5.671143e-08, 
    3.072721e-07, -4.213776e-08, 2.891186e-08, 1.917874e-08, 6.841223e-08, 
    -1.076366e-07, 5.915695e-09, -7.971664e-09, -3.025667e-09, -8.979805e-08, 
    -3.644891e-08, 8.588916e-08, 1.218191e-07, -4.207127e-08, 1.957055e-09, 
    1.955689e-08, 6.271182e-08, 1.206157e-07, 4.359429e-08, -3.348039e-08, 
    -1.660169e-09, -1.804378e-07, 1.238917e-08, -6.011042e-09, -7.208818e-08, 
    -9.047199e-10, 1.341448e-08, -1.0902e-08, 5.177345e-08, -4.538949e-08, 
    3.10456e-09, 1.228011e-08, -1.72306e-08, -3.561058e-08, 3.344007e-08, 
    -1.877299e-08, 9.9609e-09, 9.680662e-09, -2.872366e-08, 5.668344e-09, 
    3.209379e-10, 3.180196e-08, 4.071393e-08, 3.457131e-08, 1.314413e-08, 
    7.154711e-09, 1.829822e-08, 1.962377e-08, 2.630184e-07, -3.700166e-09, 
    2.193843e-07, -5.299592e-08, -6.668279e-08, -6.062908e-08, -1.30895e-07, 
    1.425428e-08, 5.127297e-08, -4.409827e-09, -3.710227e-09, 8.509232e-09, 
    -4.253396e-08, -1.031266e-07, 1.125147e-08, -6.191101e-08, -1.353267e-08, 
    -1.740398e-08, -2.099569e-09, -2.882852e-08, 6.799141e-09, 4.791787e-09, 
    -5.107142e-08, -1.119929e-09, -5.929496e-08, -2.515947e-08, 
    -5.618176e-09, -2.813181e-08, -1.428975e-08, 7.631115e-09, -1.004082e-09, 
    3.31795e-09, -1.371063e-09, 8.934634e-09, -2.340936e-09, -9.701395e-10, 
    1.11741e-07,
  -6.927089e-07, 2.397419e-07, 7.789117e-07, 1.633771e-07, -1.310768e-07, 
    -1.073204e-09, 6.452001e-08, -7.022436e-09, 6.866276e-08, -2.127672e-08, 
    3.217565e-08, 4.311255e-08, -3.522655e-08, -6.427172e-09, -2.538854e-09, 
    5.999252e-08, -9.8903e-09, 9.552878e-09, -6.896624e-08, 3.018386e-09, 
    2.233878e-08, 7.755716e-09, -1.589638e-08, 1.232047e-08, 2.611841e-08, 
    -1.602325e-08, 1.474223e-08, 1.004219e-08, -1.705985e-09, 6.377172e-08, 
    3.710784e-08, 5.452421e-10, -1.503395e-08, -2.578299e-07, -1.440117e-08, 
    6.004507e-08, -3.576424e-08, 3.161693e-08, 4.134949e-08, 6.186392e-08, 
    -7.864487e-08, 5.498396e-08, -7.927952e-09, 1.354203e-08, -4.961544e-08, 
    -4.081699e-08, 6.378843e-08, 8.124147e-08, -4.531362e-08, 1.648132e-09, 
    1.933319e-08, 4.248448e-07, 2.166723e-08, 4.400004e-08, -4.44299e-08, 
    -6.381242e-10, -1.330707e-07, -1.932131e-08, -9.453693e-09, 
    -7.689661e-08, 3.175705e-08, 5.336233e-09, -1.659491e-07, 5.795004e-08, 
    -9.666761e-08, -1.978833e-08, 2.09568e-08, -2.313391e-08, -5.032189e-08, 
    3.3986e-08, -2.54779e-08, 7.250264e-09, -7.657809e-08, -1.15399e-08, 
    2.918181e-09, 3.564537e-09, 4.044159e-08, 5.013771e-08, 2.461965e-08, 
    -3.00015e-08, 3.785442e-08, 5.394611e-09, 3.253456e-08, 4.353719e-07, 
    -2.556453e-08, 9.358064e-08, -3.523542e-08, -1.294407e-07, -5.570855e-08, 
    -1.165447e-07, 2.180514e-09, 5.129614e-08, -4.49603e-09, -1.260878e-08, 
    -4.681533e-08, -6.137869e-08, -1.325251e-07, 3.414834e-08, -5.792822e-08, 
    3.065907e-08, 6.102937e-08, -2.687553e-08, -2.928614e-08, 7.086328e-09, 
    1.742706e-08, -3.465402e-08, 5.613174e-09, -6.333357e-08, -1.690341e-08, 
    -1.006356e-09, -2.847605e-08, -1.217427e-08, 7.090421e-09, -5.818492e-10, 
    2.18165e-09, -1.601643e-09, 8.005458e-09, -2.449674e-09, -1.078575e-09, 
    -2.471916e-08,
  -4.06354e-07, 1.058875e-07, -3.869241e-08, 2.866545e-08, 1.667058e-08, 
    1.109713e-07, 6.540654e-08, 6.437176e-09, 3.784953e-08, 7.626568e-09, 
    2.19402e-08, 2.413344e-08, -4.42601e-08, 4.19891e-08, 1.645117e-08, 
    7.029523e-08, 1.892726e-09, -6.130563e-09, -3.150808e-08, 1.066496e-08, 
    1.175704e-08, 2.964953e-08, 1.935109e-08, 1.249396e-08, 2.224351e-08, 
    6.375558e-10, -1.799999e-07, 5.848051e-09, 7.679046e-08, -2.82173e-08, 
    -5.435663e-08, 3.740161e-08, -7.770154e-08, -8.868665e-08, 3.444916e-08, 
    -3.565403e-07, -3.386083e-08, 3.248121e-08, 9.119321e-08, 5.553068e-08, 
    -7.547087e-08, 3.838022e-08, -8.154245e-09, -2.802363e-09, -7.260951e-09, 
    -4.506637e-08, 7.077358e-08, 4.621972e-08, -2.959832e-08, 9.937651e-10, 
    1.925338e-08, -8.326197e-08, 1.102198e-08, 3.219666e-08, -4.725176e-08, 
    -7.089511e-10, -7.427457e-08, -3.9837e-08, -7.754739e-09, -9.183975e-08, 
    1.691546e-08, 8.499228e-10, -4.49063e-08, 3.63023e-08, -2.921452e-08, 
    1.327317e-08, 1.059902e-08, 2.20009e-08, -3.133459e-08, 4.214758e-08, 
    -2.047068e-08, 1.005219e-08, 7.702965e-09, -1.100943e-09, 3.153389e-11, 
    -2.58251e-09, 1.652657e-08, 4.383787e-08, 1.888873e-08, 7.873655e-08, 
    2.061813e-08, -6.531804e-09, 5.434083e-08, -5.155357e-08, -6.64777e-08, 
    4.151048e-08, -4.006552e-09, -1.739029e-07, -5.006826e-08, -1.122323e-07, 
    -1.543845e-08, 1.267927e-09, -3.980972e-09, 5.875085e-09, 3.392393e-08, 
    -6.367384e-08, -1.04314e-07, 4.689082e-08, -5.513743e-08, 7.694594e-08, 
    9.831388e-08, -9.224308e-09, -1.05389e-07, 7.664269e-09, -3.157129e-08, 
    -1.813873e-08, 1.086255e-08, -6.420873e-08, -3.816467e-09, 4.118192e-09, 
    -2.920615e-08, -1.094577e-08, 8.052666e-09, -4.536105e-10, 1.04933e-09, 
    -1.122544e-09, 6.880214e-09, -2.156938e-09, -1.392053e-09, -2.617594e-08,
  -1.321268e-07, 1.127603e-07, -2.257229e-08, 2.932575e-08, 5.795982e-09, 
    1.233639e-08, 2.70968e-08, 3.292621e-08, 1.805938e-08, 2.607703e-08, 
    2.917773e-08, 1.886542e-08, -5.066568e-09, 3.016157e-08, 1.889543e-08, 
    6.179789e-08, -5.522498e-09, -1.38333e-08, 4.769112e-08, 1.442481e-08, 
    8.771167e-09, 2.936258e-08, 4.107619e-08, 1.212061e-08, 2.069464e-08, 
    5.86374e-09, -1.504329e-07, 3.294053e-08, 9.876658e-09, -6.257324e-08, 
    -1.185283e-07, -1.532933e-07, 2.610909e-08, -3.465302e-07, 3.454079e-08, 
    -5.019829e-07, -3.229257e-08, 3.045488e-08, 6.107803e-08, 5.061138e-08, 
    -7.879449e-08, 2.671118e-08, -8.140262e-09, 2.067406e-09, 7.875087e-09, 
    -4.369895e-09, 5.434538e-08, 1.886974e-08, -2.919328e-08, 5.419736e-10, 
    1.946381e-08, -1.05535e-07, -2.10232e-09, 3.449736e-08, -4.644644e-08, 
    -1.843205e-09, -4.193407e-08, -5.382947e-08, -8.482672e-09, -1.18873e-07, 
    8.657253e-09, -2.651177e-10, 5.154266e-08, 3.94587e-08, 3.15913e-08, 
    1.337003e-08, -2.169622e-08, 2.291699e-08, -1.351486e-08, 5.42791e-08, 
    4.13927e-08, -9.958285e-09, 9.244332e-09, 3.740752e-09, -2.802768e-09, 
    -4.921731e-09, 2.552625e-08, 3.398253e-08, 6.571575e-09, 1.08924e-07, 
    -1.361695e-08, -1.485732e-08, 5.998038e-08, -6.598748e-08, -3.590321e-08, 
    1.239885e-07, -9.311179e-09, -1.078147e-07, -4.515374e-08, -1.232661e-07, 
    -1.954527e-08, -8.695724e-09, -5.554909e-09, 2.206323e-08, 1.041587e-07, 
    -7.664983e-08, 5.852741e-11, 1.146873e-08, -6.323626e-08, 3.808395e-08, 
    1.94294e-07, -4.905331e-09, -2.646129e-08, 8.504387e-09, -1.581302e-07, 
    -1.193712e-10, 2.393836e-08, -6.218511e-08, -3.776677e-10, 6.167056e-09, 
    -3.00131e-08, -9.847781e-09, 8.943061e-09, -1.023182e-10, 7.244125e-10, 
    -6.410119e-10, 7.830323e-09, -1.841457e-09, -1.440412e-09, -2.570414e-08,
  -2.672977e-08, 1.16919e-07, -2.048085e-08, 2.869757e-08, 8.197333e-09, 
    1.048699e-08, 9.107168e-09, 2.285839e-08, 1.228187e-08, 2.837186e-08, 
    2.380574e-08, 1.711038e-08, 1.66221e-08, 3.859651e-08, 1.989184e-08, 
    4.273602e-08, -5.386009e-08, 2.522029e-08, -1.321386e-08, 1.569055e-08, 
    7.600931e-09, 3.526731e-08, 5.070359e-08, 1.150426e-08, 1.953691e-08, 
    1.151949e-08, -1.188743e-07, 4.856969e-08, 7.613892e-09, 1.644395e-08, 
    -7.083605e-08, -4.054908e-08, -3.378562e-08, -4.427531e-07, 3.501299e-08, 
    -5.793078e-07, -3.085976e-08, 2.526146e-08, 2.885082e-08, 4.669081e-08, 
    -1.00112e-07, 2.142059e-08, -7.545538e-09, 2.775618e-09, 3.679139e-08, 
    2.221992e-08, 4.936305e-08, 5.440768e-10, -4.354286e-09, 3.308784e-10, 
    2.023754e-08, -1.112576e-07, -1.291212e-08, 3.744022e-08, -4.032088e-08, 
    -1.592014e-09, -7.451092e-09, -6.177484e-08, -9.847282e-09, 
    -9.122529e-08, 4.682704e-09, -1.39886e-09, 5.812041e-08, 6.259196e-08, 
    3.770041e-08, 1.05085e-07, -2.532789e-08, 1.099646e-07, -1.062557e-08, 
    1.949485e-08, -1.278528e-08, -1.494362e-08, 1.224106e-08, 4.830724e-09, 
    -5.487923e-09, -1.567349e-08, 2.776257e-08, 2.775488e-08, 4.473083e-09, 
    5.866019e-08, -2.782173e-08, -1.617126e-08, 6.051164e-08, -6.944884e-08, 
    2.169151e-08, -3.41409e-08, -1.016275e-08, 7.027262e-08, -4.40992e-08, 
    -1.319775e-07, -1.998109e-08, -6.35888e-09, -5.801553e-09, 2.922604e-08, 
    2.24091e-08, -8.154204e-08, 5.876235e-09, 4.74426e-08, -4.936049e-08, 
    1.627853e-08, 1.323877e-07, -3.855504e-09, -2.201074e-08, 9.377793e-09, 
    -1.279142e-07, 4.416125e-08, 2.837606e-08, -6.405759e-08, -1.93603e-09, 
    4.508536e-09, -3.049848e-08, -8.864788e-09, 1.000654e-08, 3.231548e-10, 
    -1.691831e-09, 2.269451e-09, 8.479034e-09, -1.650921e-09, -1.234113e-09, 
    -2.495136e-08,
  -1.252272e-08, 1.177665e-07, -1.945114e-08, 2.837498e-08, 7.882022e-09, 
    2.669367e-09, 6.059736e-09, 2.260583e-08, 1.048011e-08, 2.7959e-08, 
    2.191211e-08, 1.623266e-08, 2.7331e-08, 4.47136e-08, 2.004697e-08, 
    3.028269e-08, -5.254163e-08, 3.375379e-08, -2.779639e-08, 1.632759e-08, 
    6.420692e-09, 3.373657e-08, 5.226275e-08, 1.068997e-08, 1.781996e-08, 
    1.096646e-08, -9.710232e-08, 6.41686e-08, 6.730716e-09, 7.928759e-08, 
    4.224148e-09, -2.329557e-08, -3.238256e-08, -4.413664e-07, 3.530567e-08, 
    -6.320153e-07, -2.999034e-08, 1.648611e-08, 1.746571e-08, 4.369744e-08, 
    -1.039436e-07, 1.655019e-08, -6.750525e-09, 2.940755e-09, 7.49011e-08, 
    2.332888e-08, 4.461509e-08, -1.142985e-08, 2.825054e-08, -3.936051e-10, 
    2.161565e-08, -1.120912e-07, -2.274378e-08, 3.670675e-08, -2.854564e-08, 
    1.398519e-09, 9.149517e-09, -6.573778e-08, -1.143876e-08, -7.040524e-08, 
    3.196874e-09, -2.249294e-09, 6.398932e-08, 3.270918e-08, 2.191409e-08, 
    -3.56016e-08, 5.509219e-08, 8.539632e-08, -7.600761e-09, 5.785989e-08, 
    9.891096e-09, -2.17243e-08, 1.383262e-08, 4.926733e-09, -7.894197e-09, 
    -1.655565e-08, 3.181815e-08, 1.889026e-08, 1.948776e-08, -9.82925e-09, 
    -3.542448e-08, -1.773476e-08, 5.596894e-08, -7.098629e-08, 1.779529e-08, 
    -1.021606e-07, -1.01744e-08, 7.535607e-08, -4.389236e-08, -1.379798e-07, 
    -1.956244e-08, -4.940599e-10, -5.136542e-09, 2.870356e-08, -4.616095e-08, 
    -8.238045e-08, 1.60522e-08, 5.05305e-08, -3.92165e-08, 4.247319e-09, 
    1.000254e-07, -3.644637e-09, -2.922444e-08, 9.379583e-09, -5.001198e-08, 
    6.157165e-09, 2.478532e-08, -7.103142e-08, -5.029733e-09, 2.817956e-09, 
    -2.781599e-08, -7.882136e-09, 1.066212e-08, 1.053081e-09, -1.097874e-08, 
    3.50642e-09, 1.024033e-08, -1.371671e-09, -7.884324e-10, -2.381921e-08,
  -1.290545e-08, 1.176372e-07, -1.931545e-08, 2.792916e-08, 7.50066e-09, 
    9.858354e-10, 2.816876e-09, 2.197061e-08, 9.418557e-09, 2.749078e-08, 
    2.064297e-08, 1.114432e-08, 3.240422e-08, 4.769373e-08, 2.027474e-08, 
    2.801377e-08, -2.883101e-08, 4.134893e-08, -2.591135e-08, 1.674874e-08, 
    5.96566e-09, 3.219674e-08, 4.883083e-08, 1.143979e-08, 1.637653e-08, 
    1.154791e-08, -8.082083e-08, 7.537727e-08, 6.377093e-09, 1.147889e-07, 
    -3.577441e-09, 1.115035e-08, -4.044256e-08, -5.443312e-07, 3.549047e-08, 
    -6.754624e-07, -2.947047e-08, 5.541793e-09, 2.26118e-08, 4.119772e-08, 
    -1.544967e-07, 1.62002e-08, -6.086537e-09, -1.987086e-10, 7.062721e-08, 
    2.162102e-08, 4.985748e-08, -1.885348e-08, 2.479281e-08, -9.573569e-10, 
    2.323488e-08, -1.119467e-07, -2.822508e-08, 3.850295e-08, -1.801109e-08, 
    4.072831e-10, 5.243521e-09, -6.743519e-08, -1.32948e-08, -6.235646e-08, 
    2.292666e-09, -2.847798e-09, 6.744136e-08, 1.003533e-08, 1.595853e-08, 
    -2.448309e-08, 6.378656e-08, 3.850442e-08, -1.273196e-08, 8.267358e-08, 
    2.36941e-08, -2.876146e-08, 1.506788e-08, 4.522065e-09, -1.01127e-08, 
    -4.624155e-09, 3.477568e-08, 8.653359e-09, 2.409355e-08, -2.688995e-08, 
    -3.360486e-08, -1.599997e-08, 6.185832e-08, -7.199498e-08, 2.196333e-08, 
    -1.420726e-07, -9.45289e-09, 7.49904e-08, -3.495946e-08, -1.424915e-07, 
    -1.876805e-08, -5.657501e-09, -3.656623e-09, 2.3653e-08, -5.476267e-08, 
    -8.447819e-08, 2.121299e-08, 5.206795e-08, -3.145971e-08, 2.920398e-09, 
    1.044492e-07, -3.703249e-09, -3.201393e-09, 8.936091e-09, -3.160693e-08, 
    1.256393e-08, 1.793757e-08, -8.178591e-08, -9.170833e-09, 9.583232e-10, 
    -2.423457e-08, -6.313769e-09, 1.08401e-08, 1.417845e-09, -1.112784e-08, 
    1.544629e-09, 8.548014e-09, -6.404761e-10, -1.094982e-09, -2.230803e-08,
  -5.014101e-09, 1.169971e-07, -1.982238e-08, 2.737414e-08, 6.918469e-09, 
    6.86839e-10, 1.945125e-09, 2.084488e-08, 8.518043e-09, 2.687528e-08, 
    1.637585e-08, 9.048392e-09, 3.577946e-08, 4.643431e-08, 1.992834e-08, 
    4.563118e-08, -1.098085e-08, 4.392086e-08, -2.440484e-08, 1.688483e-08, 
    5.669961e-09, 3.234453e-08, 4.708846e-08, 1.141774e-08, 1.444431e-08, 
    1.144878e-08, -6.553711e-08, 5.159058e-08, 5.916661e-09, 1.348496e-07, 
    -2.267137e-08, 6.605148e-09, 4.956462e-09, -6.841076e-07, 3.578958e-08, 
    -7.083792e-07, -2.947497e-08, 3.286175e-09, 1.249481e-08, 3.971048e-08, 
    -1.573033e-07, 1.765039e-08, -5.533934e-09, -8.319407e-10, 7.047157e-08, 
    1.161646e-08, 5.69766e-08, -2.509313e-08, -7.668575e-09, -8.037944e-10, 
    2.475086e-08, -1.112265e-07, -3.076091e-08, 3.890456e-08, -1.751923e-08, 
    -1.836042e-09, 1.059055e-08, -6.790217e-08, -1.570236e-08, -5.976679e-08, 
    1.2962e-09, -3.360981e-09, 6.989995e-08, 1.880487e-09, 2.039443e-08, 
    -1.805341e-08, 8.092246e-08, 8.55801e-08, -1.594191e-08, 9.902539e-08, 
    2.691417e-08, -3.457131e-08, 1.640598e-08, 4.102219e-09, -1.23051e-08, 
    8.597851e-09, 3.568425e-08, 1.291122e-08, 2.593563e-08, -3.645033e-08, 
    -3.261505e-08, -1.551373e-08, 6.111219e-08, -7.27876e-08, 2.490953e-08, 
    -1.641341e-07, -8.476661e-09, 7.38633e-08, -2.796884e-08, -1.458761e-07, 
    -1.811071e-08, -7.717325e-09, -2.254865e-09, 1.831567e-08, -6.319084e-08, 
    -8.5642e-08, 2.522177e-08, 5.234114e-08, -2.625671e-08, 9.435901e-10, 
    1.048945e-07, -4.22088e-09, 1.54767e-08, 8.262582e-09, -1.508471e-08, 
    1.586142e-08, 4.867246e-08, -9.21537e-08, -1.355039e-08, -1.548358e-09, 
    -2.045243e-08, -3.816751e-09, 1.094048e-08, 1.642491e-09, -2.42398e-08, 
    2.432e-09, 1.2301e-08, -2.459117e-09, -4.678569e-09, -2.134453e-08,
  -4.98909e-09, 1.157908e-07, -1.911172e-08, 2.665882e-08, 6.465427e-09, 
    9.723067e-10, 2.07109e-09, 1.934637e-08, 7.64129e-09, 2.580697e-08, 
    1.250822e-08, 1.268694e-08, 3.758504e-08, 4.445332e-08, 1.964401e-08, 
    5.403763e-08, -9.745236e-09, 4.464482e-08, -2.301027e-08, 1.646043e-08, 
    5.382219e-09, 3.202337e-08, 4.682983e-08, 1.090308e-08, 1.315829e-08, 
    1.113182e-08, -5.739793e-08, 4.514487e-08, 5.532399e-09, 1.464225e-07, 
    -4.410941e-08, 9.587382e-09, 2.388009e-08, -7.490819e-07, 3.642145e-08, 
    -7.334965e-07, -3.012861e-08, 4.106013e-09, 4.535707e-09, 3.874974e-08, 
    -1.445532e-07, 1.900077e-08, -5.03772e-09, -4.848154e-09, 7.904117e-08, 
    1.206837e-08, 5.74322e-08, -2.92751e-08, -3.521724e-08, -2.243887e-09, 
    2.651146e-08, -1.09914e-07, -3.142245e-08, 4.017014e-08, -2.54992e-08, 
    -3.514799e-09, 2.363134e-08, -6.778372e-08, -1.903625e-08, -5.781312e-08, 
    -3.166178e-11, -3.289813e-09, 7.108252e-08, 7.557894e-09, 2.232683e-08, 
    -1.724351e-08, 8.334854e-08, 1.022842e-07, -1.797031e-08, 1.132058e-07, 
    4.319571e-08, -1.000427e-08, 1.74303e-08, 3.717957e-09, -1.458474e-08, 
    2.622556e-08, 3.523034e-08, 1.446278e-08, 2.414687e-08, -3.976646e-08, 
    -3.36733e-08, -1.544542e-08, 5.453177e-08, -7.330999e-08, 2.261669e-08, 
    -1.739779e-07, -7.695974e-09, 7.199657e-08, -2.101348e-08, -1.486096e-07, 
    -1.736004e-08, -5.183245e-09, -1.087471e-09, 1.370207e-08, -6.713714e-08, 
    -8.614383e-08, 2.739463e-08, 5.178953e-08, -2.29316e-08, 6.801066e-10, 
    1.035503e-07, -4.667143e-09, 1.554001e-08, 7.41084e-09, -1.680235e-09, 
    1.886923e-08, 2.143938e-07, -9.89566e-08, -1.661573e-08, -5.488062e-09, 
    -1.835264e-08, -1.113278e-09, 1.093525e-08, 1.779824e-09, -5.189219e-08, 
    8.663733e-10, 1.077879e-08, -8.219203e-11, -4.632788e-09, -1.987263e-08,
  -4.771323e-09, 1.135812e-07, -2.000752e-08, 2.522279e-08, 5.865331e-09, 
    1.313083e-09, 2.910724e-09, 1.705882e-08, 6.488904e-09, 2.44828e-08, 
    1.076069e-08, 1.363458e-08, 3.696573e-08, 4.372146e-08, 1.906142e-08, 
    6.397406e-08, -8.950394e-09, 4.459281e-08, -2.155097e-08, 1.653871e-08, 
    4.952653e-09, 3.116713e-08, 4.614253e-08, 9.976702e-09, 1.17567e-08, 
    1.008755e-08, -5.440313e-08, 4.125513e-08, 5.134666e-09, 1.565854e-07, 
    -4.741605e-08, 4.793378e-09, 2.967829e-08, -8.944852e-07, 3.752928e-08, 
    -7.504527e-07, -3.131148e-08, 3.287568e-09, -7.92727e-09, 4.296652e-08, 
    -1.296887e-07, 1.995693e-08, -4.584422e-09, -3.456108e-09, 8.278676e-08, 
    1.36971e-08, 5.764184e-08, -3.259635e-08, -4.398785e-08, -2.888207e-09, 
    2.933416e-08, -1.076463e-07, -3.091776e-08, 4.032445e-08, -3.048468e-08, 
    -8.951417e-09, 2.568174e-08, -6.860235e-08, -2.431398e-08, -5.716085e-08, 
    -1.832746e-09, -2.631964e-09, 7.09872e-08, -1.817639e-10, 2.35329e-08, 
    -1.589558e-08, 8.125846e-08, 1.229594e-07, -1.181854e-08, 1.27214e-07, 
    5.439483e-08, -3.279922e-08, 1.822139e-08, 3.470973e-09, -1.744947e-08, 
    -1.773981e-08, 3.701892e-08, 1.65083e-08, 2.188578e-08, -4.090441e-08, 
    -3.689416e-08, -1.511281e-08, 4.664781e-08, -7.359199e-08, 2.265517e-08, 
    -1.772016e-07, -6.415803e-09, 6.895357e-08, 4.98607e-09, -1.522178e-07, 
    -1.613625e-08, -3.905643e-09, -3.077787e-10, 9.56967e-09, -6.904372e-08, 
    -8.538515e-08, 2.339302e-08, 5.043296e-08, -2.008994e-08, 4.041567e-10, 
    1.025356e-07, -4.934037e-09, 1.024246e-08, 6.518505e-09, 1.324997e-08, 
    2.264892e-08, 1.370364e-07, -1.022488e-07, -1.8234e-08, -8.770485e-09, 
    -1.917363e-08, -2.582965e-10, 1.172305e-08, 1.318995e-09, -6.3377e-08, 
    7.407835e-11, 1.052041e-08, 4.848388e-10, 1.32149e-08, -1.760725e-08,
  -4.101366e-09, 1.083923e-07, -2.39047e-08, 2.205309e-08, 4.55816e-09, 
    1.938815e-09, 5.493348e-09, 1.189017e-08, 4.116259e-09, 2.198271e-08, 
    8.727852e-09, 1.191052e-08, 3.406035e-08, 4.114509e-08, 1.759827e-08, 
    5.811108e-08, -7.085146e-09, 4.340689e-08, -1.918382e-08, 1.702278e-08, 
    3.955961e-09, 2.866238e-08, 4.458366e-08, 8.090524e-09, 9.045038e-09, 
    7.296194e-09, -4.548292e-08, 3.803609e-08, 4.57112e-09, 1.552215e-07, 
    -4.773335e-08, -3.703235e-09, 3.132595e-08, -9.593944e-07, 4.017988e-08, 
    -7.457515e-07, -3.284858e-08, 4.92723e-09, -1.637966e-08, 4.446085e-08, 
    -1.096897e-07, 1.997091e-08, -4.219146e-09, -3.090388e-09, 8.084726e-08, 
    1.747492e-08, 6.369726e-08, -3.526594e-08, -4.236344e-08, -1.272102e-08, 
    3.290012e-08, -1.025609e-07, -2.93418e-08, 3.974519e-08, -2.110411e-08, 
    -2.188523e-08, 1.938247e-09, -6.963841e-08, -3.546703e-08, -5.740016e-08, 
    -5.174002e-09, -1.14585e-09, 6.959863e-08, -1.502119e-08, 3.087801e-08, 
    -1.339174e-08, 8.097436e-08, 1.191956e-07, -1.114813e-08, 1.340677e-07, 
    5.984839e-08, -9.262703e-08, 1.908245e-08, 2.861725e-09, -2.291103e-08, 
    9.339374e-10, 3.262593e-08, 1.638477e-08, 2.251266e-08, -3.986474e-08, 
    -2.278631e-08, -1.450754e-08, 4.166861e-08, -7.322751e-08, 2.555032e-08, 
    -1.778143e-07, -3.700734e-09, 6.237451e-08, -7.744184e-09, -1.44406e-07, 
    -1.281126e-08, -3.912351e-09, -2.618208e-10, 6.591131e-09, -6.966798e-08, 
    -8.210323e-08, 3.263538e-08, 4.690094e-08, -1.726437e-08, 3.446772e-10, 
    1.048661e-07, -5.051341e-09, 4.318295e-09, 5.65943e-09, 1.437343e-08, 
    2.985814e-08, 1.012371e-07, -1.037184e-07, -1.886315e-08, -1.013325e-08, 
    -1.95887e-08, 1.671197e-11, 9.497171e-09, 1.72588e-09, -6.542314e-08, 
    -5.081915e-10, 1.040459e-08, -1.131878e-08, 1.113371e-08, -1.341903e-08,
  1.337341e-13, 9.008071e-14, 1.412175e-13, 2.317488e-13, 3.243202e-13, 
    4.068268e-13, 1.850706e-13, -2.242523e-13, -3.758736e-13, 1.25671e-12, 
    3.900744e-13, -1.203613e-14, -3.607825e-13, 4.348487e-13, 2.629433e-14, 
    -3.608527e-14, 6.669967e-13, -1.331964e-13, -2.097704e-13, -8.629045e-13, 
    -3.017317e-12, -5.572171e-13, 6.003418e-13, -1.082523e-12, 4.587366e-14, 
    1.426505e-13, 6.750328e-14, 5.584879e-14, 4.140353e-14, -1.662063e-13, 
    -1.256505e-14, -1.837626e-13, -1.503906e-13, -1.88697e-13, -1.951139e-13, 
    -4.249896e-13, 9.22948e-13, -2.245409e-12, 2.454872e-14, -3.416308e-13, 
    1.403169e-12, -1.637815e-14, -2.437631e-13, -6.250012e-15, 2.599716e-13, 
    4.216571e-13, -3.765349e-14, 8.421334e-13, -9.09654e-13, 1.256554e-12, 
    5.959481e-13, -2.66444e-15, 4.732901e-13, -1.083766e-12, -2.233681e-13, 
    -2.35525e-12, -1.141079e-13, -4.030667e-13, 3.247894e-13, 1.555196e-12, 
    9.033398e-13, -2.684076e-13, 3.334171e-13, 7.834938e-13, 1.750827e-13, 
    -5.604692e-13, -1.360687e-13, 2.090442e-13, -1.637544e-13, 1.802299e-13, 
    -1.13353e-13, 4.005029e-14, -1.280018e-13, -1.097104e-13, -6.285164e-13, 
    -5.876712e-13, 2.407427e-13, 2.062864e-15, 7.205672e-14, -1.931755e-13, 
    -1.908725e-12, 5.603329e-13, -1.366751e-13, -1.571313e-14, 1.583734e-13, 
    2.399367e-15, -9.348145e-13, 4.034216e-13, -4.476649e-13, 3.051276e-13, 
    -6.174891e-14, 5.910379e-13, -1.903412e-13, -7.281725e-14, -1.227609e-13, 
    -2.865064e-13, -3.430854e-14, 1.002489e-13, -2.762661e-14, -9.690796e-13, 
    3.57981e-13, -7.2021e-14, -7.447338e-13, 9.301598e-13, 1.065577e-13, 
    5.064487e-13, 6.821332e-13, 2.976524e-13, 3.876855e-13, 2.437239e-13, 
    1.971727e-13, 7.873103e-15, -5.330819e-15, 2.373473e-14, 3.915362e-13, 
    -3.218895e-12, -8.403022e-13, -7.785193e-13, -2.205234e-12, 7.233283e-14,
  -3.973237e-13, -3.829181e-13, -2.841532e-13, -2.046614e-13, -2.103798e-13, 
    -2.433862e-13, -2.330815e-13, -1.28085e-13, -3.426112e-13, 1.323069e-14, 
    -2.446656e-13, 2.068284e-14, 4.835431e-13, 4.772463e-13, 5.035557e-13, 
    2.072538e-13, -1.20775e-13, -4.267787e-13, -2.292945e-13, -5.373148e-13, 
    -7.163134e-13, -6.90571e-13, -3.36776e-13, -8.812463e-16, -2.352879e-14, 
    -1.033027e-13, -3.012027e-13, -3.548935e-14, 1.358063e-14, -1.17312e-13, 
    -3.340776e-13, -1.05688e-13, 2.232833e-13, -1.092214e-13, -7.682354e-14, 
    -3.120409e-14, 1.143251e-12, 2.196791e-13, -8.956488e-14, -6.00963e-13, 
    -2.008059e-12, -1.076825e-13, -3.17779e-13, -7.791982e-14, 4.092722e-13, 
    3.107572e-13, -1.863672e-12, 6.516251e-13, 3.121622e-13, 9.466385e-13, 
    -2.993494e-13, -2.730163e-15, 3.938879e-13, 8.011695e-13, 3.097368e-14, 
    -3.143045e-13, 9.595361e-14, -1.837376e-12, -1.246236e-12, 3.830077e-12, 
    6.491738e-13, -3.794596e-13, 5.057321e-14, -1.927469e-13, -3.773653e-13, 
    -5.972467e-14, -3.915978e-13, -1.083401e-14, 5.629765e-13, 5.586463e-13, 
    9.252856e-13, -2.161587e-13, 1.950496e-13, 2.508233e-13, -1.216223e-12, 
    -1.497623e-12, 5.287763e-13, 5.776527e-13, -5.55465e-13, -2.372951e-13, 
    -8.647305e-13, -3.443664e-13, 6.286233e-13, -2.134029e-13, -3.292525e-13, 
    -4.770782e-13, 7.186002e-13, 3.538607e-13, -3.400795e-13, 8.024927e-14, 
    -2.80498e-13, -1.59462e-12, 1.094507e-12, -8.500777e-13, -7.917948e-14, 
    1.162692e-13, -4.795888e-13, 5.448389e-13, 2.705013e-13, -6.469803e-13, 
    -2.259667e-13, 5.615868e-13, 4.636475e-13, -5.900557e-12, -1.982872e-13, 
    -7.515106e-13, -2.64006e-13, -1.895984e-12, -1.355274e-12, -3.037367e-13, 
    4.663051e-14, 1.718457e-13, 1.415141e-13, -3.808075e-14, 1.582905e-13, 
    -5.386151e-13, -4.807935e-12, 4.270204e-13, 2.953067e-14, 1.653551e-14,
  6.77236e-15, 9.582612e-14, 8.778395e-14, 1.03445e-13, 6.344231e-14, 
    -6.664808e-14, -2.621028e-13, -2.364081e-13, -1.582762e-14, 
    -9.145462e-14, 1.854072e-14, 1.660963e-13, -1.70676e-13, -1.623007e-13, 
    1.288553e-14, 5.185602e-13, 1.644296e-13, 1.037018e-13, 4.249309e-13, 
    8.809203e-13, 4.688541e-13, 3.850253e-13, 9.25468e-13, 4.270612e-13, 
    6.315781e-13, 5.489845e-13, -3.213402e-13, 6.886852e-14, 1.581721e-13, 
    3.002251e-13, -1.473127e-14, -1.125627e-13, -2.913156e-13, -1.991671e-13, 
    8.400919e-14, 7.042283e-14, 6.21625e-13, 3.582083e-13, -1.763173e-14, 
    -9.776367e-13, 1.853817e-12, 2.278039e-14, -2.381845e-13, 3.500796e-13, 
    -5.516212e-13, 1.953299e-14, -6.517946e-13, -2.10813e-12, 1.012579e-13, 
    1.709262e-13, -4.536441e-13, 3.677683e-13, -1.421761e-12, -6.157677e-12, 
    2.98675e-13, 1.689579e-12, 1.060693e-12, -1.435421e-13, -7.761604e-13, 
    -5.01931e-13, -5.071915e-13, -9.00377e-13, 1.502479e-13, 2.880598e-13, 
    2.228093e-13, 1.584705e-13, -4.406198e-14, 6.188106e-14, -5.89806e-14, 
    -3.404568e-13, 1.972755e-12, 1.650763e-14, -1.12306e-12, 1.68178e-13, 
    -4.759381e-13, -1.288476e-12, -6.443205e-13, 1.02484e-13, 1.328697e-11, 
    1.952188e-13, 9.302975e-14, 6.070161e-14, -1.059718e-12, 6.109557e-13, 
    3.387499e-13, -1.880926e-13, 8.76646e-13, 9.067053e-13, -3.449176e-13, 
    -2.086602e-12, -1.034173e-13, -3.165093e-13, 3.418307e-13, -2.885049e-12, 
    8.820028e-14, -4.369886e-13, -8.690618e-13, 2.954581e-13, 1.00437e-12, 
    7.06862e-12, -1.132136e-12, -3.299323e-13, 6.35633e-13, -1.714062e-12, 
    6.347006e-14, 5.60274e-13, 1.05644e-12, 2.053309e-12, 2.196611e-12, 
    1.804869e-12, 1.193358e-12, 5.892994e-13, 4.287334e-13, 1.324635e-14, 
    5.000098e-13, 2.533593e-12, 3.702724e-13, 1.593513e-12, -1.827101e-12, 
    -1.766087e-13,
  7.452372e-15, 1.584011e-13, 8.511247e-14, -1.533496e-13, -3.341355e-13, 
    -3.849698e-13, -2.908507e-13, -8.626433e-14, -1.165734e-15, 9.894863e-14, 
    2.328276e-13, -3.319983e-13, -2.023659e-13, 3.961553e-13, 3.240186e-13, 
    2.484443e-13, 1.13104e-14, 6.938894e-15, 4.88054e-13, -1.292438e-13, 
    -1.013495e-13, 8.921197e-13, 1.566081e-12, 1.130901e-13, -6.701584e-14, 
    -6.794565e-14, 4.621303e-15, -1.068867e-13, 1.903477e-13, -2.416123e-14, 
    9.258427e-13, 3.308603e-13, 8.14071e-14, -3.162748e-14, 3.188977e-13, 
    1.61246e-13, -1.116707e-12, 1.49384e-13, 9.391099e-14, -1.537509e-12, 
    1.0696e-12, 2.74919e-13, -2.962283e-13, 3.067754e-13, 2.435413e-13, 
    -6.294965e-14, -6.841749e-15, -1.292355e-12, -3.885503e-13, 
    -1.483754e-12, -1.170904e-13, -1.318737e-12, -1.492263e-12, -4.07524e-12, 
    9.071407e-13, 2.388902e-12, -4.153719e-12, 3.335887e-13, 3.282555e-13, 
    -1.928699e-12, -8.995443e-13, -7.457368e-13, -2.714495e-14, 4.789502e-14, 
    2.702283e-14, -3.865241e-13, -9.896112e-13, -6.33868e-13, -6.815937e-13, 
    -4.073408e-13, 1.302333e-12, 1.126182e-13, 6.15244e-13, -9.10938e-14, 
    -1.382333e-12, -2.849249e-13, 1.946672e-13, 1.379553e-12, 3.298033e-12, 
    3.917699e-14, 3.636536e-13, -2.517754e-12, 3.428924e-13, 6.104006e-13, 
    9.794943e-14, -3.079897e-13, -6.555728e-13, -1.040223e-12, -1.070442e-12, 
    -1.484063e-12, -3.781281e-13, 2.643441e-13, 3.535228e-13, 8.512011e-13, 
    -9.411916e-14, -1.163378e-11, -1.102865e-12, -1.713768e-13, 4.583833e-13, 
    -7.776002e-13, -8.948536e-13, -8.942456e-13, 4.164741e-13, -6.112697e-13, 
    2.603473e-14, 3.476247e-13, 5.755951e-13, 7.848583e-13, 7.975842e-13, 
    5.026535e-13, 8.552742e-13, 4.785061e-13, 2.699369e-13, -6.826484e-14, 
    -4.922035e-13, 3.095962e-12, -7.383504e-12, 3.533207e-13, -2.915003e-13, 
    1.133815e-13,
  -1.182665e-13, -1.546124e-13, -1.539047e-14, -9.056644e-14, -1.821876e-13, 
    -1.781908e-13, -3.097383e-13, -4.420908e-13, -1.489087e-13, 1.88341e-12, 
    5.855733e-13, 8.03288e-13, 1.765532e-13, 1.179612e-13, -3.503725e-13, 
    1.428885e-13, -1.981609e-14, -4.537343e-13, -1.549993e-13, -2.63678e-13, 
    -1.246586e-12, -4.363176e-14, 9.741097e-13, 4.11185e-13, 4.431316e-13, 
    2.163131e-13, 5.915129e-13, -3.219786e-13, -5.143108e-14, 6.059042e-14, 
    3.54633e-13, 1.219622e-12, 2.366579e-13, 3.070461e-13, -1.659964e-12, 
    -4.882622e-13, -6.448425e-13, -3.63997e-13, 5.003914e-13, -1.160976e-12, 
    -2.546824e-13, -2.020883e-12, 1.42171e-13, -4.043554e-13, 4.710177e-12, 
    -1.394287e-12, -2.029904e-13, -1.372558e-12, -5.817957e-13, 5.421944e-12, 
    1.976128e-13, -2.671988e-12, -1.13842e-12, 3.369804e-13, 8.20434e-13, 
    4.533408e-12, -1.653733e-12, 1.489822e-13, -1.861927e-13, -2.118965e-14, 
    -9.651169e-13, -4.558992e-13, -4.433537e-13, -1.061484e-13, 
    -7.145951e-14, -5.573181e-13, -2.366163e-13, -3.312767e-13, 
    -3.373829e-13, -2.769035e-13, 8.003181e-13, -3.558265e-14, -1.900147e-13, 
    -3.177875e-13, -1.58096e-12, -8.469336e-13, -4.578837e-13, -4.272971e-13, 
    1.551832e-12, -6.106227e-16, 1.104512e-12, 5.103265e-13, 7.911727e-14, 
    -2.429085e-12, -6.095124e-13, 1.655995e-12, -1.183359e-12, 4.193867e-14, 
    -1.168439e-12, -1.616041e-12, -4.516665e-13, 1.817754e-12, 3.307493e-13, 
    6.761355e-13, -2.795125e-13, 3.068176e-12, -1.848383e-13, 3.164968e-13, 
    2.977188e-12, -1.879386e-13, -1.199554e-12, -2.061741e-12, 2.505617e-13, 
    5.79049e-13, -4.070494e-13, 5.640488e-13, 5.157819e-13, 4.793943e-13, 
    8.432144e-13, 3.783085e-13, 8.118506e-15, 4.205802e-13, 1.631612e-13, 
    6.84855e-13, -1.48323e-12, 2.704682e-12, 2.530564e-12, -6.501149e-12, 
    -2.030866e-12, -5.062756e-13,
  -2.918221e-13, -4.418133e-13, -4.11754e-13, -4.326539e-13, -3.285705e-13, 
    -3.925749e-13, 2.214617e-13, -2.796374e-13, 2.087414e-12, 9.096057e-13, 
    -2.87298e-13, -1.647016e-13, 2.944034e-13, 1.163986e-12, 3.463729e-12, 
    2.027573e-13, 1.290273e-13, -2.564476e-13, -1.185586e-12, -1.184969e-12, 
    -1.187883e-12, 1.10445e-12, 2.563588e-12, 9.48075e-13, -5.878631e-13, 
    -1.01183e-12, 7.251422e-13, -5.967449e-15, 5.791478e-13, -1.409706e-12, 
    -9.604539e-13, 2.791933e-12, 2.767037e-12, 1.068173e-12, -3.341216e-13, 
    2.438882e-13, 1.81255e-13, -2.281439e-13, -8.847645e-13, -8.402251e-13, 
    7.347012e-13, -1.285758e-11, -2.672862e-13, -7.333392e-13, 1.362538e-11, 
    1.62817e-12, -7.270573e-14, -4.195463e-13, 7.939371e-13, 1.413389e-11, 
    1.077929e-12, -4.988315e-12, -4.753448e-13, -7.340017e-12, 6.445511e-13, 
    4.30217e-12, 4.006795e-13, -3.424788e-13, -6.724537e-13, 4.824353e-12, 
    1.754236e-12, -5.042661e-12, -2.045863e-13, -1.636469e-14, 2.676137e-13, 
    1.936229e-13, -1.847134e-13, -4.083872e-12, -2.081946e-12, 5.900752e-12, 
    7.04381e-13, 5.61412e-13, -6.01158e-13, -1.445066e-12, -2.433337e-12, 
    -9.055257e-13, -1.30819e-13, -1.014966e-12, -1.47087e-12, -2.412709e-12, 
    1.647266e-12, 1.066774e-12, 6.893514e-13, -1.440154e-12, 1.147721e-12, 
    3.510664e-12, 6.759537e-12, -2.411682e-13, -1.172572e-12, -7.126244e-13, 
    8.421042e-14, 1.259676e-12, 3.308326e-13, -3.059092e-12, 1.599221e-12, 
    5.564271e-13, -1.248807e-12, -4.235778e-13, 1.823122e-11, 9.970635e-13, 
    1.55273e-12, 4.016718e-13, 1.035536e-12, 4.529556e-12, -9.340306e-13, 
    -4.513889e-13, -1.582068e-15, 3.525236e-13, -9.603429e-15, 4.96464e-13, 
    -9.539591e-14, 4.254097e-13, 4.833633e-13, 2.151085e-12, -1.544181e-12, 
    1.506131e-12, 1.037307e-11, -1.158745e-11, -1.041105e-12, -3.027301e-12,
  1.691425e-13, 2.566281e-13, 3.939071e-13, 7.654988e-13, 3.946843e-14, 
    -2.651768e-13, 2.871592e-12, -4.8761e-13, 1.742773e-12, 1.904199e-12, 
    4.40592e-13, -3.448519e-12, 4.862277e-12, 4.872103e-12, 1.014117e-11, 
    -2.105149e-13, 9.204914e-13, -1.335015e-12, -2.086553e-12, -1.266875e-12, 
    -1.953993e-13, 1.626477e-14, 1.292855e-13, 6.47038e-13, -2.639e-12, 
    -4.964584e-12, 8.797962e-13, -7.989664e-12, -5.323519e-14, -4.310829e-12, 
    -1.289246e-11, -3.839928e-12, 3.511968e-12, -5.045242e-12, -1.154299e-12, 
    -2.193357e-12, 4.92717e-13, -2.700895e-13, 1.761868e-12, -1.665279e-13, 
    -3.804157e-12, -9.077405e-12, -9.432871e-13, -1.055723e-12, 3.049783e-12, 
    -1.399214e-12, -7.653322e-13, -8.690826e-13, 2.358669e-13, 1.230303e-11, 
    9.954745e-13, -1.437128e-12, -5.318135e-13, -5.069001e-12, 7.928047e-13, 
    2.694234e-13, 2.197575e-12, -5.247469e-14, -1.381489e-12, 1.763895e-12, 
    -5.713208e-13, 1.813993e-12, 1.722456e-12, 1.38467e-12, 9.38838e-13, 
    7.345236e-13, -4.475365e-12, 3.685274e-12, 1.404266e-12, 1.083689e-11, 
    -2.105538e-13, 4.747314e-13, 1.899592e-13, -1.007305e-12, -2.623135e-12, 
    -3.106959e-13, 3.646458e-13, -1.974615e-12, -1.727132e-12, -4.419742e-12, 
    -9.691914e-12, -2.214237e-12, 9.399426e-13, -9.168777e-13, 5.318523e-13, 
    4.028333e-12, 7.253642e-12, 4.795608e-13, -4.015798e-14, -9.598711e-13, 
    2.659151e-12, -4.098499e-12, 2.518818e-14, -5.189382e-12, -3.847644e-12, 
    -7.258083e-14, -1.346445e-12, -2.036704e-12, 2.602585e-12, 2.399969e-13, 
    5.333123e-12, 1.659402e-12, 6.218463e-13, 4.938758e-13, 4.712897e-14, 
    -3.924638e-13, -3.759215e-13, -1.470157e-12, -1.163958e-12, 1.532108e-14, 
    -1.047384e-12, -1.059763e-12, -5.265621e-12, -3.916978e-12, 
    -6.095457e-12, 3.539491e-12, 9.345372e-12, 5.411895e-12, 1.880093e-14, 
    2.773892e-12,
  2.017608e-12, 2.824962e-12, 2.600975e-12, 2.305489e-12, -3.018641e-12, 
    -8.175127e-12, -3.581746e-12, 2.154338e-11, 1.567252e-11, 1.938161e-11, 
    3.49436e-11, 3.050232e-11, 2.096112e-11, 1.840644e-11, 5.727974e-12, 
    -9.410251e-14, -5.101936e-12, -9.253709e-14, -9.646867e-13, 
    -1.387779e-12, 2.405298e-13, 1.471545e-12, 4.944378e-13, -6.913359e-13, 
    7.984169e-13, 3.542999e-12, -3.638201e-12, -5.324075e-13, 3.466116e-12, 
    -5.846601e-12, -1.27609e-11, 5.74929e-13, -3.997802e-12, -9.25926e-12, 
    -4.584721e-12, -1.506295e-12, 2.822675e-12, -5.955861e-13, 2.689454e-11, 
    -5.910994e-13, -4.918055e-12, -1.89726e-12, 3.765988e-12, 7.68516e-12, 
    -2.051304e-12, 2.211675e-12, -2.110701e-12, -4.085066e-13, 5.681089e-12, 
    1.069987e-11, -6.511874e-13, 8.066381e-12, -5.83078e-13, 7.542211e-12, 
    2.256029e-13, -5.259126e-13, 1.140094e-11, -7.284507e-13, -2.411343e-12, 
    -3.895342e-12, -9.510726e-13, 4.970357e-12, 4.281575e-12, -3.295708e-12, 
    -3.01803e-12, -8.932355e-12, -1.670963e-11, 1.034367e-11, 5.043799e-12, 
    -1.334322e-12, -5.487e-12, -3.011924e-12, 3.943401e-12, -8.01248e-12, 
    -1.361594e-12, 2.663425e-13, 4.023934e-13, -1.84823e-12, -1.687001e-12, 
    -9.277579e-12, -4.268083e-11, 1.063343e-11, -2.82574e-12, 3.421985e-12, 
    4.646838e-13, 1.28399e-11, 2.007949e-12, -3.038236e-12, -8.439898e-13, 
    -4.350964e-13, 1.082745e-12, 6.633916e-12, 1.965234e-13, -2.412071e-13, 
    -1.184719e-12, 3.21399e-12, -2.305378e-12, -3.336276e-12, -1.815936e-12, 
    -2.695732e-13, 1.33904e-12, 2.136378e-12, -3.240186e-13, -8.097793e-13, 
    -4.243828e-13, -6.988854e-13, -1.110778e-13, -3.65924e-12, -6.18372e-12, 
    -9.235945e-13, -6.848133e-12, -8.180345e-12, -1.392458e-11, 
    -3.769096e-12, -4.408696e-12, 1.708724e-11, 9.465428e-12, -1.770363e-12, 
    4.750367e-14, 1.430628e-11,
  2.106454e-12, 7.556705e-12, 1.192912e-11, -1.906808e-14, -4.536677e-12, 
    2.516723e-11, 3.966177e-11, -9.171552e-13, -2.138134e-11, -7.935763e-12, 
    1.425851e-11, 8.341244e-12, -7.099876e-14, 7.141399e-12, -4.916345e-13, 
    -9.201675e-12, -7.012807e-13, -3.775036e-13, 2.385203e-12, 4.519524e-12, 
    3.948647e-12, 4.55655e-12, 6.361328e-12, 9.569651e-12, 1.239464e-11, 
    2.690828e-11, 6.993156e-12, -5.365697e-11, -7.761042e-12, -2.563483e-11, 
    -2.300968e-11, 1.332748e-11, 1.892153e-12, 6.470102e-13, 2.614881e-12, 
    4.488687e-12, 2.206471e-12, -2.54758e-13, 1.385975e-11, -4.686113e-13, 
    2.576028e-12, -3.98237e-13, 6.356922e-12, 9.287805e-13, -1.377376e-11, 
    9.379442e-12, 3.554185e-12, -1.440001e-12, 8.053814e-12, 1.583907e-11, 
    -1.774223e-12, -3.60989e-13, -1.743272e-12, 9.475487e-12, -2.307578e-13, 
    -8.479328e-14, 3.359507e-12, -3.13774e-13, 1.693473e-12, -8.140173e-12, 
    2.617268e-12, 6.741413e-12, -4.883566e-12, 1.225353e-13, 2.497891e-13, 
    6.304457e-12, -5.14852e-12, 3.954226e-12, 2.674458e-11, -5.614539e-11, 
    -1.334155e-12, 1.789291e-12, 9.557632e-13, -1.235309e-11, 1.462919e-12, 
    2.234324e-14, 7.22547e-14, -3.244588e-11, -2.61458e-12, 6.110668e-12, 
    -3.79982e-11, 4.732139e-12, -2.555497e-12, 1.922651e-11, 1.31864e-12, 
    1.395564e-11, -2.170125e-12, -1.873338e-11, -3.539452e-13, -3.553546e-13, 
    4.91085e-12, -8.923196e-13, 6.744952e-13, -2.275402e-13, -8.925305e-12, 
    -3.740841e-13, -2.595701e-13, -7.046308e-12, -9.350576e-13, 
    -1.187533e-12, -1.622985e-11, -1.8658e-11, 1.606874e-13, -3.334572e-12, 
    -6.115997e-12, 1.225603e-12, 3.864131e-13, 5.048267e-12, -4.162337e-12, 
    -5.856843e-12, -4.266421e-12, -6.852657e-12, 6.043221e-12, 7.758461e-12, 
    7.836232e-13, 2.373913e-11, 6.962004e-12, -1.514394e-12, -6.494666e-13, 
    7.910478e-12,
  3.595414e-11, -4.786602e-12, -3.27248e-12, -9.109616e-12, 1.864216e-11, 
    7.035129e-11, -7.279552e-12, -3.769766e-11, -2.147089e-11, -2.726612e-11, 
    1.482499e-11, -6.734488e-12, 8.79348e-12, 7.130893e-12, 7.266146e-12, 
    -8.460913e-12, -1.650879e-12, 4.837075e-12, 4.894241e-12, 6.575199e-12, 
    4.457837e-12, 5.441134e-12, 1.272825e-11, 1.654968e-12, 6.983455e-12, 
    -4.375181e-12, 1.536153e-11, -9.391224e-12, 1.003199e-11, -1.310184e-11, 
    -2.216256e-11, -2.486525e-12, 1.879039e-12, 1.387987e-12, 1.326038e-11, 
    2.058492e-13, -4.73982e-13, 4.438533e-13, -1.621604e-11, -1.249059e-12, 
    1.529207e-12, -1.24846e-12, 7.673737e-12, -1.194903e-12, 4.560755e-12, 
    1.506226e-12, 5.157111e-12, 1.064315e-12, 3.005388e-12, 1.261757e-11, 
    -2.243056e-12, 1.704761e-12, -2.55328e-12, 1.10407e-12, -9.830664e-13, 
    1.516287e-13, -3.586839e-12, 1.26015e-12, 3.294012e-12, -4.871045e-12, 
    -9.303044e-12, 2.877185e-12, 9.405671e-13, -1.565118e-12, 1.638514e-12, 
    -3.378173e-12, -7.675235e-12, 1.219512e-11, 8.766335e-12, 2.737828e-11, 
    -3.770456e-13, -3.954753e-13, 1.596209e-12, 1.277851e-11, 5.290809e-12, 
    6.415701e-14, -1.016201e-13, 1.182027e-12, -2.654459e-12, 1.33767e-11, 
    -2.537565e-11, -1.833414e-12, 3.236383e-12, -6.101605e-12, -1.708005e-11, 
    4.068204e-12, 1.061998e-12, -2.602406e-11, 5.478504e-13, 1.811051e-14, 
    2.651587e-12, -7.049083e-14, 1.387758e-12, 1.594344e-12, -1.283459e-12, 
    5.243042e-12, 7.489481e-13, 1.945104e-11, 5.222031e-12, -4.43752e-12, 
    -2.310499e-12, -1.531449e-11, 1.260556e-12, -4.442401e-12, 1.630376e-12, 
    1.433451e-12, 6.881509e-12, 8.015325e-12, 5.629316e-12, -1.258375e-11, 
    4.58171e-12, -3.74957e-12, 1.18499e-11, 7.298676e-12, -4.058934e-12, 
    1.013612e-11, 3.117836e-12, -1.543874e-12, 2.971035e-12, 4.994796e-12,
  1.005057e-10, -6.15748e-11, -4.310585e-11, -4.575895e-12, 3.995876e-11, 
    9.37983e-12, -4.289824e-11, -3.518547e-11, 4.241246e-11, 3.748724e-12, 
    -1.64696e-12, -1.609873e-11, -2.358053e-11, 7.871481e-14, 7.141343e-12, 
    -2.569772e-12, -5.120626e-13, 8.213957e-12, 5.691489e-12, 3.108569e-12, 
    2.271239e-12, 7.16488e-12, 1.372708e-11, 1.972089e-12, -1.661171e-12, 
    -2.081813e-11, -5.646705e-12, -2.541051e-11, 2.823852e-12, 2.898615e-11, 
    -8.584627e-11, -2.197614e-11, -3.404443e-12, 3.997858e-12, 2.143519e-11, 
    9.192092e-12, -7.71927e-13, 9.545767e-13, -1.324897e-10, 5.404566e-14, 
    -2.39353e-13, -7.368828e-12, -1.771222e-13, -7.995939e-13, 8.484546e-12, 
    -7.035539e-12, 4.247186e-12, 1.99013e-12, 2.866707e-13, 3.535335e-12, 
    -1.287902e-11, 3.072292e-11, 7.036482e-13, 2.860601e-13, 1.773109e-12, 
    2.705336e-13, -2.087391e-11, 2.247985e-12, 6.535983e-12, -1.252044e-11, 
    -1.681422e-11, -2.158662e-12, 1.215805e-12, 1.547418e-12, 5.045564e-12, 
    -1.286193e-13, -1.8825e-11, 3.796241e-12, -2.48932e-11, 5.637363e-11, 
    1.759998e-11, -9.450385e-12, 2.47341e-12, -8.159806e-12, 1.408723e-12, 
    6.000755e-14, 3.146233e-13, 2.80741e-11, -1.0623e-12, 5.738132e-12, 
    -1.524922e-11, 3.419487e-14, 4.551193e-12, -3.305634e-11, -2.668143e-12, 
    -2.006578e-11, 4.625023e-12, -8.554379e-12, 4.800145e-13, -9.504619e-13, 
    2.880474e-13, 9.011791e-12, 7.50372e-14, 7.796081e-12, 2.099526e-11, 
    9.132745e-12, 1.074695e-14, 1.592043e-11, 3.207046e-12, -6.192224e-12, 
    1.332201e-11, -3.202751e-13, 1.459211e-12, -2.192364e-12, 1.176353e-11, 
    2.63044e-11, 3.182987e-11, 2.242434e-11, 8.511802e-12, -9.364731e-12, 
    8.762713e-12, 1.307487e-11, 3.371248e-12, 1.966149e-12, -5.270007e-12, 
    -2.128464e-13, 8.466075e-13, -1.708291e-12, 5.275523e-12, -2.243183e-11,
  1.709255e-11, -6.702816e-11, -4.745626e-11, -5.524914e-12, -2.227307e-11, 
    -4.970535e-11, -4.589551e-11, -3.416822e-11, 1.552203e-11, 1.649192e-11, 
    -3.149658e-11, -9.633561e-11, -1.158318e-11, -6.110956e-11, 
    -5.920375e-12, -3.767342e-12, -3.368306e-12, 1.030087e-11, 3.383377e-12, 
    -6.161072e-12, -5.471845e-12, 1.110712e-11, 1.095501e-11, 5.385692e-12, 
    1.057732e-11, -2.872969e-11, 4.337863e-12, 2.672773e-11, 1.148837e-11, 
    -1.862954e-11, 4.080158e-11, -4.188361e-11, -3.080958e-11, 3.013412e-11, 
    7.342948e-11, -2.811507e-11, 1.158496e-12, 1.080247e-13, -3.620961e-10, 
    1.17375e-12, 8.51319e-13, -1.455924e-11, -6.724121e-12, -4.72327e-13, 
    -9.170664e-12, 1.170242e-11, 3.267386e-12, 6.762368e-13, 1.247891e-14, 
    1.737915e-13, -2.100306e-11, 2.209988e-11, 2.726375e-12, 1.751221e-12, 
    1.342115e-12, 2.493561e-13, -2.12943e-11, 4.376055e-13, 3.325873e-12, 
    -2.331524e-12, -7.993606e-13, 5.595524e-14, 1.867284e-11, 8.716139e-13, 
    8.745316e-12, -3.822986e-11, -1.863176e-11, -5.503709e-11, 1.602496e-12, 
    2.69671e-11, -6.043077e-11, -1.567828e-10, -2.872835e-11, 7.114309e-13, 
    -3.198708e-12, 2.597922e-14, 6.278034e-13, 1.573253e-11, 2.730427e-13, 
    -3.71192e-12, -1.070888e-11, 5.862422e-13, -1.898037e-12, -2.384137e-11, 
    1.675993e-11, 5.242229e-11, 1.280687e-11, 8.812062e-12, -7.993294e-13, 
    -2.626344e-12, 1.742295e-11, 1.615552e-11, -8.194001e-13, 1.344893e-11, 
    1.25564e-11, 9.81224e-12, -3.506528e-13, -3.454126e-12, 1.942224e-12, 
    -3.370149e-12, 1.203837e-11, 6.858333e-12, 1.476319e-12, -3.535228e-13, 
    5.385559e-11, 6.947132e-11, 6.017764e-11, 4.216894e-11, 2.454259e-12, 
    -1.503708e-11, 5.968115e-12, 2.533262e-11, 5.187406e-12, 1.968425e-12, 
    1.215406e-11, -4.739986e-13, 6.444845e-14, -1.124691e-12, 2.915487e-12, 
    9.666046e-12,
  -6.063683e-11, -5.334555e-11, -6.846079e-11, -5.370326e-11, -5.195622e-11, 
    -4.866796e-11, -2.67264e-11, 1.698908e-11, 2.253622e-10, 3.60707e-11, 
    -9.571743e-11, -1.663292e-10, 1.779887e-11, -5.480283e-12, -9.905321e-11, 
    -6.608847e-12, 3.926948e-12, 6.716294e-12, -4.006295e-12, -1.125122e-11, 
    -7.024381e-12, 8.598011e-12, 6.773027e-12, 3.863243e-11, -5.431233e-11, 
    -1.275091e-11, 2.45497e-11, 9.224399e-12, 2.072986e-11, 3.092171e-11, 
    3.760903e-11, -5.975531e-11, -1.729945e-10, -2.504241e-11, 1.041065e-10, 
    7.226042e-11, 3.01803e-13, -2.409184e-14, -2.599425e-10, 5.193845e-13, 
    -4.794654e-12, -2.036971e-11, -1.231559e-11, 2.58106e-13, -7.753576e-11, 
    5.340461e-11, 1.824874e-12, 8.399392e-13, 9.072743e-14, 8.537615e-14, 
    -2.957287e-11, 8.045298e-11, 5.416556e-13, 2.354517e-12, -4.489409e-13, 
    1.64091e-13, -1.470837e-10, -7.293499e-13, -2.292815e-11, 1.364531e-11, 
    3.419331e-11, 1.932343e-11, 3.137668e-11, 1.579359e-11, 2.178124e-11, 
    -7.629763e-11, -1.069078e-11, -9.357359e-11, -2.335931e-11, 
    -4.103606e-11, -8.432699e-11, -1.693325e-10, 1.112215e-10, -2.734812e-11, 
    -2.372058e-12, 3.796963e-14, 7.234491e-13, 5.890899e-12, 6.291579e-13, 
    3.008038e-12, -7.655321e-12, -7.288825e-12, -5.908496e-12, -3.83622e-11, 
    5.154543e-12, 1.363252e-10, -3.754175e-11, 1.853317e-11, -2.290473e-12, 
    -2.274181e-12, 2.185674e-11, 1.711675e-11, -6.135648e-13, 2.034324e-11, 
    -5.859313e-12, 8.36069e-12, -2.074696e-12, -6.796785e-11, 5.795142e-12, 
    -1.759259e-12, -1.729283e-11, 2.622409e-11, 7.929629e-13, 8.167078e-14, 
    7.522138e-11, 1.284128e-10, 1.277316e-10, 5.872725e-11, -1.366462e-11, 
    -2.352851e-11, 8.419709e-12, 3.635492e-11, 9.523493e-12, 4.568568e-12, 
    2.482659e-11, -2.78888e-14, -1.26732e-13, -3.039236e-13, 6.571965e-13, 
    4.376366e-11,
  -6.796919e-11, -7.093304e-11, -9.381518e-11, -5.914513e-11, -3.113776e-11, 
    -2.878808e-11, 5.464962e-12, 1.715086e-10, 3.909175e-10, 2.120393e-11, 
    -1.25171e-10, -1.785132e-10, 3.510969e-11, 4.532197e-11, -3.191949e-10, 
    -4.846523e-12, 1.432094e-11, 1.500888e-11, -2.167871e-11, -1.521228e-11, 
    -1.048539e-11, 4.298784e-12, 1.060574e-11, 1.945955e-11, -1.025491e-11, 
    -1.11255e-10, 3.980594e-11, -1.805889e-11, 1.460121e-11, -6.051915e-11, 
    1.033484e-10, -9.046053e-11, -1.737721e-10, 2.471001e-11, 2.342522e-10, 
    2.019718e-10, -1.894707e-12, 2.28928e-13, -1.342189e-10, 8.542944e-13, 
    -2.284031e-11, -2.393952e-11, -1.375633e-11, -4.060155e-13, 
    -2.652834e-10, 5.227863e-11, -4.136691e-13, 4.015899e-12, -2.729372e-13, 
    6.681322e-13, -1.295375e-11, 7.076073e-11, 8.548273e-12, 4.35767e-12, 
    -3.283373e-13, 1.64313e-14, -2.100395e-10, 4.511058e-13, -4.463106e-11, 
    3.883671e-12, 6.947065e-11, 3.950618e-11, 1.439515e-11, 2.180283e-11, 
    1.630811e-11, -1.342131e-10, 5.341061e-12, -1.763536e-10, -5.035217e-11, 
    6.052048e-12, -1.099694e-10, -7.809975e-11, -3.108314e-11, -1.299858e-10, 
    3.305001e-12, -1.558753e-13, 3.247957e-13, -3.58602e-14, 5.255685e-13, 
    1.728706e-11, -6.430856e-12, -7.692213e-12, -6.329159e-12, -2.286531e-10, 
    -1.857403e-11, -1.720433e-10, -1.57327e-10, 2.859091e-11, -1.38313e-12, 
    -1.490807e-12, 7.469092e-11, 5.144596e-12, -1.979528e-13, 1.571334e-11, 
    -3.39222e-11, 3.776535e-12, -5.439649e-12, -1.37315e-10, 1.559908e-11, 
    -9.998224e-13, -7.152057e-11, 5.952011e-11, 1.466605e-13, -2.640665e-13, 
    6.75775e-11, 2.056093e-10, 2.502802e-10, 9.652679e-11, -9.84457e-12, 
    -2.333111e-11, 1.541789e-11, 4.026246e-11, 1.216582e-11, 1.015321e-11, 
    1.988054e-11, 1.138201e-13, 6.500356e-14, 1.104394e-13, -4.828637e-13, 
    3.08451e-11,
  -7.181478e-11, -1.116158e-10, -1.244811e-10, -5.941314e-11, -2.772116e-11, 
    6.017187e-12, 9.114287e-11, 2.872651e-10, 5.028411e-10, -3.377587e-11, 
    -1.597897e-10, -1.326603e-10, -1.433742e-12, 7.138001e-11, -2.551472e-10, 
    5.21494e-13, 1.433826e-11, 1.292455e-11, -3.48459e-11, -1.58773e-11, 
    -8.874013e-12, 2.892575e-12, 8.04401e-12, -9.997447e-11, 2.150347e-11, 
    1.411198e-10, 9.330092e-12, 1.404721e-11, 8.172019e-11, -2.025269e-12, 
    2.888931e-10, -8.333623e-11, -2.988145e-10, 1.616287e-10, 5.106766e-10, 
    4.437826e-10, -3.874456e-12, 3.667067e-13, -2.132323e-10, 1.051381e-12, 
    -4.121934e-11, -8.395284e-12, -7.305712e-12, -1.923336e-12, 
    -5.949323e-10, 1.003442e-11, -5.175638e-12, 2.813971e-12, 9.236611e-13, 
    1.577127e-12, 3.230971e-11, 6.283396e-11, 2.907394e-11, 8.397683e-12, 
    2.345901e-13, -6.150636e-14, -6.045142e-11, 6.41962e-12, -4.955001e-11, 
    -2.972877e-11, 8.638668e-11, 4.56768e-12, 1.882827e-11, 2.038365e-11, 
    2.693716e-11, -1.228229e-10, -1.467761e-10, -3.432385e-10, -1.08803e-10, 
    -5.761813e-11, -6.371814e-11, -1.908875e-10, 1.027334e-11, -1.109257e-10, 
    1.004481e-11, -4.363176e-13, -9.969803e-14, -1.262479e-11, -3.752288e-12, 
    -4.809331e-11, -5.771605e-12, 1.01692e-12, -5.391021e-12, -5.106877e-10, 
    -3.475908e-11, -3.466116e-13, -2.134315e-11, 3.574008e-11, -3.401446e-13, 
    -2.542633e-12, 1.343243e-10, 9.761391e-12, 3.641532e-14, 1.139138e-11, 
    -4.399081e-11, -6.262324e-12, -1.046385e-11, 2.031928e-10, 2.016853e-11, 
    -8.734791e-13, -1.175142e-10, -6.805895e-11, -9.80882e-14, -8.667511e-13, 
    1.024671e-10, 2.71698e-10, 4.730258e-10, 1.523863e-10, -1.899036e-11, 
    -1.335398e-11, 2.653944e-11, 3.86986e-11, 8.685275e-12, 1.255507e-11, 
    8.21454e-12, -7.092105e-14, -6.816769e-14, -2.262635e-13, -1.588174e-12, 
    1.17788e-11,
  -7.967471e-11, -1.448732e-10, -1.219413e-10, -5.732015e-11, 4.827472e-12, 
    7.590484e-11, 8.288148e-11, 2.858205e-10, 5.252752e-10, -8.432166e-11, 
    -2.857596e-10, -1.070144e-11, -8.562551e-11, 1.516942e-11, 8.43301e-11, 
    2.144729e-12, 1.08201e-11, -3.253176e-12, -3.65622e-11, -5.828893e-12, 
    1.121103e-12, 4.72089e-12, -1.491918e-12, -1.483487e-10, -1.262768e-12, 
    1.539464e-10, 5.850276e-11, 1.381146e-10, 1.237412e-10, -1.377856e-10, 
    4.671874e-10, 1.769476e-10, -2.534433e-10, 4.507055e-10, 3.491014e-10, 
    3.318477e-10, -6.446621e-12, 3.860245e-13, -5.003089e-10, -2.952971e-12, 
    -3.801381e-11, 2.94762e-11, 6.803003e-12, -2.931252e-12, -8.165839e-10, 
    4.017453e-12, -2.142508e-12, -1.188716e-11, 5.963985e-12, 3.381739e-12, 
    9.390277e-11, 1.107126e-10, 4.605974e-11, 1.436313e-11, -4.237277e-13, 
    1.800782e-13, 1.255416e-10, 1.959122e-11, -4.157256e-11, -1.630113e-10, 
    9.117174e-11, -5.013745e-11, -1.226093e-10, 3.962559e-11, 4.256137e-11, 
    2.004319e-10, -2.91507e-10, -2.589482e-10, -1.873965e-10, -5.187117e-11, 
    4.877454e-11, -1.271536e-09, 1.698306e-10, -8.583134e-12, 2.240559e-11, 
    -1.419975e-12, -1.660894e-13, -2.278866e-11, -1.364195e-11, -1.51976e-10, 
    -6.756595e-12, 4.725664e-12, 1.063816e-12, -8.153662e-10, -1.652392e-10, 
    -4.566727e-10, -1.953582e-10, 3.948153e-11, 1.006834e-13, -6.907586e-12, 
    1.048026e-10, 5.449938e-11, 3.752332e-12, 1.159917e-12, 3.838196e-11, 
    -5.979439e-12, -1.720468e-11, 3.172549e-10, 1.945488e-11, -4.32876e-12, 
    -5.68503e-11, -1.51084e-10, -4.687917e-13, -2.144063e-12, 1.056544e-10, 
    5.284664e-10, 8.830165e-10, 4.531808e-10, -1.28686e-11, -9.043211e-12, 
    4.014855e-11, 3.028799e-11, 3.202993e-12, 6.589618e-12, 8.528511e-12, 
    4.751754e-15, 6.328271e-14, -8.049672e-13, -3.444134e-12, -8.362e-11,
  -9.015366e-11, -1.888765e-10, -1.569411e-10, -8.275869e-11, 4.099121e-11, 
    1.029719e-10, 1.35465e-11, 2.072849e-10, 4.443894e-10, 9.993251e-11, 
    -7.434533e-10, -8.742163e-11, -1.725429e-10, -1.462688e-10, 
    -1.710099e-10, 7.532463e-12, 3.855227e-12, -5.581313e-12, -2.600764e-11, 
    1.157652e-11, 1.470646e-11, 5.25624e-12, -4.174439e-13, -1.807088e-11, 
    -1.689262e-10, -1.816733e-10, 4.459331e-10, -1.380798e-10, 3.346301e-10, 
    3.106226e-10, 9.137313e-10, 5.974439e-10, -1.434959e-10, 4.055529e-10, 
    2.710188e-10, 3.235812e-10, -7.609913e-12, 4.0834e-13, -8.866543e-10, 
    -1.708429e-11, 1.066134e-11, 6.716938e-11, 2.112355e-11, 1.516315e-12, 
    -7.03329e-10, 1.140599e-11, 1.605027e-11, -2.260681e-11, 1.030607e-11, 
    6.876499e-12, 2.099338e-10, -2.225153e-10, 1.010836e-10, 2.36998e-11, 
    -1.025269e-12, 2.158274e-13, 8.039791e-11, 4.275034e-11, -3.804441e-11, 
    -4.390424e-10, 8.757617e-11, -3.95417e-12, -3.305072e-10, 5.620002e-11, 
    2.838121e-11, 1.633715e-10, -4.714131e-10, -9.775469e-11, -3.553247e-10, 
    1.823253e-11, 1.272937e-11, -2.395005e-09, -5.787548e-11, 8.459011e-12, 
    8.99993e-11, -3.112177e-12, 1.74083e-13, -2.797806e-11, -1.990679e-11, 
    -2.246932e-10, -9.372947e-12, 1.923128e-12, 2.05409e-11, -7.752945e-10, 
    -4.934098e-10, -9.620322e-10, -1.120029e-10, 2.620659e-11, 6.198653e-13, 
    -1.53122e-11, -7.486811e-11, 6.254304e-11, 1.265699e-11, 3.995755e-11, 
    1.75989e-10, 1.018918e-11, -2.519407e-11, 2.097504e-10, 1.343636e-11, 
    -1.255884e-11, 1.469598e-10, -1.708835e-10, -2.317702e-12, -5.324963e-12, 
    1.4386e-10, 6.35227e-10, 1.192584e-09, 1.073584e-09, 7.704415e-11, 
    -7.078782e-12, 6.060574e-11, 1.972644e-11, -1.941913e-11, -1.838352e-11, 
    4.172485e-11, 3.355538e-13, 3.587131e-12, -9.829915e-13, -5.208722e-12, 
    -2.978933e-10,
  -8.311041e-11, -2.252758e-10, -3.221441e-10, -1.943299e-10, 5.160672e-11, 
    7.477396e-11, -1.476685e-11, 4.908607e-11, 3.023128e-10, 7.248424e-11, 
    -1.092159e-09, -1.64512e-10, -2.277964e-10, -2.85107e-10, -4.55687e-10, 
    1.821707e-11, -5.656453e-12, 2.726708e-11, -6.527223e-12, 2.103029e-11, 
    2.794565e-11, 6.53344e-12, 1.975486e-11, 1.603429e-10, -3.414744e-10, 
    -8.514007e-10, 8.74147e-10, -1.427566e-09, -2.57927e-11, -4.695799e-11, 
    2.437643e-09, 2.96545e-10, -3.223217e-10, 8.954331e-10, 1.040315e-09, 
    3.587211e-10, -1.024425e-12, -4.218847e-14, -9.742482e-10, -4.189094e-11, 
    -5.237162e-11, 6.985346e-11, 2.125011e-11, 2.010192e-11, -7.255032e-10, 
    3.557687e-11, 5.856293e-11, -2.492762e-11, 8.776269e-12, 1.437173e-11, 
    3.007039e-11, -8.680932e-10, 2.643677e-10, 3.798881e-11, 8.408385e-13, 
    -3.552714e-14, 3.677769e-11, 7.562306e-11, -6.946674e-11, -4.736509e-10, 
    7.674572e-11, 2.12232e-10, -3.310205e-10, 4.900329e-11, 1.464571e-11, 
    1.574207e-10, -5.461303e-10, -8.447465e-11, -6.784777e-10, -4.29619e-10, 
    -1.731024e-10, -2.552323e-09, -5.182912e-10, -2.193481e-10, 5.652703e-10, 
    -8.597567e-13, 6.96776e-13, -1.205258e-11, -1.880647e-11, -2.589999e-10, 
    -1.835065e-11, -2.398348e-12, 5.167777e-11, -7.485816e-10, -5.7865e-10, 
    -1.749214e-10, 1.196785e-10, 2.532019e-11, 1.288941e-12, -4.154188e-11, 
    -1.93781e-10, 3.636274e-11, 2.148903e-11, 2.726575e-10, 1.696563e-10, 
    2.965095e-11, -3.534062e-11, 1.268656e-10, 6.068035e-12, -2.766321e-11, 
    2.704148e-10, -6.391565e-11, -4.852341e-12, -1.26078e-11, 2.625935e-10, 
    3.031619e-10, 8.315872e-10, 1.74019e-09, 2.883329e-10, 5.488943e-13, 
    8.049739e-11, 5.547562e-12, -4.837553e-11, -4.517275e-11, 1.224709e-10, 
    9.784173e-13, 1.389333e-11, -8.98781e-13, -5.134004e-12, -3.268124e-10,
  3.311662e-10, -2.934151e-10, -4.203855e-10, -3.966321e-10, -4.090595e-11, 
    3.832312e-11, 2.887646e-11, -9.534773e-11, 3.194458e-10, -2.471054e-10, 
    -1.008189e-09, -3.632898e-10, -2.604565e-10, -4.32486e-10, -7.407728e-10, 
    3.729603e-11, -2.594334e-11, 6.427747e-11, 1.188738e-11, 1.870148e-11, 
    3.653255e-11, 1.722356e-11, 5.751843e-11, 2.183853e-10, -4.542322e-10, 
    -1.698336e-09, 9.183907e-10, -1.263814e-09, 1.183658e-10, 3.672888e-09, 
    1.914007e-09, 7.0618e-10, -1.283105e-09, 1.633701e-09, 1.853056e-09, 
    4.583924e-10, -8.512302e-13, -2.614797e-12, -1.0081e-09, -7.38332e-11, 
    -7.030323e-11, 3.756995e-11, 8.808954e-12, 6.000139e-11, -1.552536e-09, 
    8.829915e-11, 3.137988e-10, -5.191403e-12, -3.171152e-12, 3.10485e-11, 
    -7.971401e-13, -8.575327e-10, 4.79303e-10, 5.024461e-11, -9.089529e-12, 
    3.801404e-13, -2.605667e-10, 1.039833e-10, -1.365862e-10, -2.801266e-10, 
    7.035439e-11, 2.999663e-10, -1.292442e-10, 3.277378e-11, 5.370282e-12, 
    -1.64043e-10, -2.879261e-10, 2.672707e-11, -1.031243e-09, -8.118626e-10, 
    -5.367617e-10, -1.722753e-09, 2.775593e-10, -3.74353e-10, 2.030907e-09, 
    8.835599e-12, 1.101785e-12, -7.042367e-12, -2.621796e-11, -2.406466e-10, 
    -5.156764e-11, -1.209193e-11, 9.485568e-11, -6.398295e-10, 6.339107e-11, 
    -8.9031e-12, 2.18769e-10, 5.650236e-11, 8.142376e-13, -1.060982e-10, 
    -3.368932e-10, 2.189452e-10, 2.517186e-11, 6.52263e-10, 4.100329e-10, 
    2.163176e-11, -4.573479e-11, 3.698091e-10, -5.091039e-12, -8.687807e-12, 
    4.411902e-10, -3.978595e-11, -4.583667e-12, -2.374478e-11, 3.48539e-10, 
    2.87983e-11, 3.373515e-10, 2.215657e-09, 4.747385e-10, 2.358647e-11, 
    1.002363e-10, -1.76712e-11, -1.101803e-10, -6.022915e-11, 2.340883e-10, 
    2.136602e-12, 3.637313e-11, 1.009193e-13, -2.310596e-12, -3.178258e-11,
  5.621139e-10, 3.247855e-10, 1.115161e-10, -2.035669e-10, -2.549818e-10, 
    -1.535838e-11, 8.50271e-11, -4.172769e-10, 4.769198e-10, -3.702461e-10, 
    -4.483276e-10, -5.048513e-10, -2.550173e-10, -7.041372e-10, 
    -1.128274e-09, 4.814851e-11, -1.067093e-11, 7.892353e-11, 2.008971e-11, 
    2.170708e-12, 3.05711e-11, 2.470202e-11, 6.874856e-11, 2.06807e-10, 
    -2.495391e-10, -2.860549e-09, 9.640324e-10, 6.604601e-10, 2.448648e-09, 
    4.774162e-09, 4.955645e-10, 1.700482e-09, -2.781544e-09, 1.787893e-09, 
    1.83088e-09, 4.193232e-10, -3.805312e-11, -5.594636e-12, -3.043713e-09, 
    -2.291479e-10, 1.321048e-10, -6.663115e-11, -6.558309e-12, 1.241455e-10, 
    -6.467253e-10, 2.036948e-10, 1.831587e-09, 1.926708e-10, -1.450289e-11, 
    6.83249e-11, -1.914255e-10, 9.424888e-10, 7.144543e-10, 4.160867e-11, 
    -5.460201e-11, 1.367795e-12, 4.035563e-10, 1.172893e-10, 6.748472e-10, 
    -3.910747e-10, 6.813039e-11, 1.808367e-10, -5.216059e-10, 1.908163e-11, 
    1.753833e-11, -8.474466e-10, 1.700009e-10, -3.775504e-10, -9.608421e-10, 
    -2.910053e-09, -9.772272e-10, -8.124594e-10, -2.711609e-10, 
    -2.700808e-10, 2.853553e-09, 1.66942e-11, 1.071143e-12, -3.231548e-11, 
    -5.532481e-11, -2.144809e-10, -1.342073e-10, -1.68038e-11, 1.39714e-10, 
    -1.601457e-10, -8.268231e-11, 5.13932e-10, -5.848833e-11, 1.140954e-10, 
    -3.647305e-12, -1.975451e-10, -7.303846e-10, 5.941935e-10, 2.020073e-11, 
    8.74423e-10, 9.690027e-11, -3.756355e-11, -5.290062e-11, 8.035279e-10, 
    -2.210854e-11, 5.242597e-11, 2.211742e-10, -1.00564e-11, -1.058709e-12, 
    -3.479972e-11, 5.555059e-10, 3.393907e-11, -9.465495e-11, 1.615728e-09, 
    5.424639e-11, -2.026717e-10, 1.043823e-10, -3.914735e-11, -2.183818e-10, 
    -1.014406e-10, 3.606964e-10, 4.237677e-12, 6.876455e-11, 2.576384e-12, 
    3.126388e-13, 2.73122e-10,
  6.233698e-10, 4.768488e-10, 7.29937e-10, 7.121592e-10, 2.189999e-10, 
    1.00151e-11, 5.670486e-11, -6.525518e-10, 6.871623e-10, -1.138805e-09, 
    -1.305953e-09, -8.228973e-10, -1.589378e-10, -9.795862e-10, -1.65377e-09, 
    -3.014833e-11, 2.923883e-12, 1.346194e-10, 1.005951e-11, -3.373302e-11, 
    1.651657e-11, 2.227907e-11, 6.462031e-11, 1.798206e-10, 9.908128e-10, 
    -4.267665e-09, 2.380904e-09, 7.671979e-10, 2.304642e-09, 3.170275e-09, 
    2.092296e-09, 3.092349e-09, -2.295256e-09, 2.054332e-09, 1.888043e-09, 
    1.623295e-09, -1.803585e-10, -2.948752e-12, -9.00776e-09, -5.027389e-10, 
    4.268692e-10, -2.760565e-10, -2.281197e-11, 2.119449e-10, 2.215014e-09, 
    3.97943e-10, 4.236913e-09, -4.911271e-11, -1.072991e-11, 7.325918e-11, 
    -1.998295e-10, 2.601038e-09, 6.078154e-10, -2.637179e-11, -1.273881e-10, 
    1.392664e-12, 3.135234e-10, 1.830095e-10, -4.545356e-10, -2.709784e-09, 
    3.821654e-11, 5.084999e-11, -3.503651e-10, 2.381952e-11, 3.378986e-11, 
    -1.161499e-09, -8.806147e-10, -1.885265e-09, -1.026525e-09, -1.85381e-09, 
    -8.136887e-10, 6.136709e-10, 4.017444e-10, 3.954277e-10, 2.018034e-09, 
    8.878231e-12, 1.231015e-12, -2.213518e-11, -7.723368e-11, -2.601546e-10, 
    -2.772396e-10, -1.084253e-11, 1.30715e-10, -2.485226e-09, 1.177476e-10, 
    6.199876e-10, -6.177636e-10, 1.501839e-10, -2.731815e-12, -2.706884e-10, 
    -1.288623e-09, 6.482375e-10, 1.659117e-12, 8.566218e-10, -5.564367e-10, 
    -1.116433e-10, -7.07935e-11, 6.681624e-10, -5.601564e-11, 1.300371e-10, 
    6.831833e-10, 1.919389e-10, 6.221246e-12, -4.773559e-11, -4.911378e-10, 
    2.883418e-10, -2.16108e-10, 2.630784e-11, 1.377725e-09, -1.359194e-09, 
    9.702816e-11, -2.762235e-11, -3.665939e-10, -2.503207e-10, 4.979235e-10, 
    4.563816e-12, 6.706902e-11, 3.938849e-12, -3.648637e-12, 2.197673e-10,
  6.242118e-10, 1.507203e-10, 1.855966e-09, 1.113563e-09, 1.020069e-09, 
    6.217249e-10, 3.809646e-10, -2.526122e-10, 8.748628e-10, -2.274192e-09, 
    -1.619313e-09, 1.091635e-09, -5.550618e-10, -4.370264e-10, -1.990387e-09, 
    -2.457398e-10, 2.472689e-11, 3.435545e-10, 2.401634e-12, -7.416645e-11, 
    2.113154e-11, 3.012701e-11, 4.617107e-11, 6.346568e-11, 8.933227e-10, 
    -5.243706e-09, -1.416851e-09, -2.045965e-09, 1.151534e-09, 1.493859e-09, 
    4.133227e-09, 4.213945e-09, -1.130417e-09, 2.29241e-09, 1.8631e-09, 
    2.155318e-09, -3.165681e-10, 4.563461e-12, 2.541924e-09, -3.815799e-10, 
    9.60793e-10, -3.913669e-10, -5.641709e-11, 3.201202e-10, 6.812883e-09, 
    6.622685e-10, 4.27773e-09, 9.841017e-11, -4.115464e-12, 1.583711e-11, 
    -9.501733e-11, 1.507132e-09, 2.088583e-10, -1.854289e-10, -2.043308e-10, 
    -2.40874e-12, 2.59206e-11, 5.192845e-10, -1.567254e-09, -3.562683e-09, 
    -4.092726e-12, 1.291767e-11, 1.749072e-09, 4.087326e-11, 8.690222e-11, 
    -1.327308e-09, 2.963532e-10, 3.118117e-09, -3.373898e-09, -2.438114e-09, 
    -6.828031e-10, 1.170079e-09, 3.269491e-10, 3.24124e-09, 1.133213e-09, 
    -2.839329e-11, 2.67697e-12, 6.927436e-11, 2.382627e-11, -7.76339e-11, 
    -4.625988e-10, -3.979182e-11, -1.504219e-11, -1.227541e-08, 
    -1.926992e-10, -1.164452e-09, -6.991598e-10, 1.686118e-10, 4.652367e-11, 
    -1.884217e-10, -1.120597e-09, 7.582115e-10, -2.249934e-11, 6.89667e-10, 
    -1.259963e-09, -1.661306e-10, -1.265221e-10, -1.738698e-10, 
    -1.154206e-10, 1.70715e-10, 1.473026e-09, 6.276668e-10, 1.370548e-11, 
    -7.402257e-11, 4.359777e-09, 6.552625e-10, 1.885496e-10, 8.464411e-10, 
    -8.482459e-10, -2.111022e-10, -1.04535e-10, -1.196554e-11, -6.55902e-10, 
    -6.455707e-10, 6.383658e-10, -5.334755e-12, -5.073808e-11, -3.521627e-12, 
    -2.599698e-11, 2.403056e-11,
  8.151027e-10, -8.963532e-10, 3.389584e-09, 9.085106e-10, 1.266582e-09, 
    1.268898e-09, 1.530122e-09, 1.28173e-09, 1.6211e-09, -1.771912e-09, 
    -3.313634e-09, 5.152824e-09, -3.887841e-10, 1.577572e-09, -2.237559e-09, 
    -4.005379e-10, 9.131682e-11, 6.766747e-10, 6.984102e-11, -8.592238e-11, 
    4.49738e-11, 1.486846e-10, 4.451906e-11, 4.335412e-10, -1.858712e-09, 
    -7.251106e-09, -9.517613e-10, -5.184123e-09, 7.57634e-10, 5.441869e-10, 
    1.48424e-08, 8.443347e-09, 4.789591e-10, 1.796106e-09, 1.799545e-09, 
    4.163905e-09, 3.038778e-11, 1.35163e-11, 4.131703e-09, -5.722639e-11, 
    1.738641e-09, -2.954756e-10, 3.719691e-11, 4.32449e-10, 9.169067e-09, 
    9.844108e-10, 4.777601e-09, -1.532037e-10, -2.874359e-11, -1.802656e-10, 
    4.603802e-10, 2.383693e-10, 1.593399e-10, -1.171685e-12, -3.538553e-10, 
    -9.34719e-12, -9.413448e-10, 1.950575e-09, 3.190202e-10, 4.604228e-10, 
    -6.014744e-12, -3.14806e-11, -7.719692e-11, -2.401073e-10, 1.710156e-10, 
    -2.735437e-09, 6.537526e-10, -1.210143e-09, -4.773842e-09, -2.971351e-09, 
    3.309673e-10, 4.867182e-10, 2.541292e-10, 3.217988e-09, 2.871575e-09, 
    -8.884982e-11, 4.646949e-12, 1.560814e-10, 1.397837e-10, 1.205745e-09, 
    -6.623075e-10, -1.400647e-10, -2.325571e-10, -2.751148e-08, 
    -1.544638e-09, 1.454563e-09, -2.275335e-10, 1.712515e-10, 2.205325e-10, 
    2.173017e-10, -2.000924e-10, 9.214935e-10, -1.548273e-11, 8.065946e-10, 
    -2.160679e-09, -2.036579e-10, -2.240974e-10, -8.44711e-10, -2.001777e-10, 
    1.958306e-10, 1.135472e-09, 1.154524e-09, 1.568878e-11, -1.121849e-10, 
    1.078123e-08, 4.284395e-10, 6.186376e-10, 1.684295e-09, -6.270433e-10, 
    -3.174836e-09, -9.780372e-10, 1.080984e-10, -1.077797e-09, -9.339693e-10, 
    8.412648e-10, 1.939782e-13, -7.987921e-11, -2.872147e-11, -4.108891e-11, 
    7.318235e-11,
  1.722498e-09, -2.253273e-09, -2.781348e-10, -1.024119e-09, -3.794298e-11, 
    1.76658e-09, 2.908564e-09, 3.073495e-09, 3.330399e-09, 2.966488e-09, 
    -1.739522e-09, 1.212129e-09, 2.605418e-10, 7.133849e-11, -2.410189e-09, 
    -7.315009e-10, -1.156451e-10, 1.186706e-09, 2.028955e-11, -5.647394e-11, 
    1.162448e-11, 4.418723e-10, 9.742962e-11, -6.66688e-10, -3.37684e-09, 
    -1.177287e-08, -2.66067e-09, -6.710906e-09, -4.925766e-10, -1.878334e-09, 
    2.496233e-08, 1.532015e-08, -2.291245e-09, 1.916817e-09, 7.561312e-10, 
    7.413149e-09, 3.629509e-10, 2.646416e-11, 6.297398e-09, -9.094435e-10, 
    3.003987e-09, -7.784706e-11, 4.466258e-10, 6.965504e-10, 6.748394e-09, 
    1.126665e-09, -7.171366e-09, -1.255863e-09, -1.350998e-10, -2.351985e-10, 
    5.062191e-10, 8.714096e-11, 3.269264e-10, -6.408527e-11, -4.567404e-10, 
    -1.377032e-11, -2.494403e-09, 5.070075e-09, -6.256192e-09, 2.360245e-10, 
    1.813305e-11, -1.247713e-10, -2.704894e-10, -1.227193e-09, 1.894193e-10, 
    -4.574872e-09, 6.400569e-11, -3.669072e-09, -1.03872e-08, -3.670579e-09, 
    9.280541e-10, -1.827033e-09, -8.506618e-11, 3.586933e-09, 6.995938e-09, 
    -1.69706e-10, 1.383427e-11, 2.21128e-10, 1.010292e-10, 1.736765e-09, 
    -8.516849e-10, -3.192355e-10, -2.564633e-10, -2.14695e-08, 1.296598e-10, 
    5.7139e-10, 1.04572e-09, 1.494129e-10, 6.225025e-10, 5.994565e-10, 
    8.472512e-11, 1.593969e-09, 3.402789e-11, 1.222264e-09, -3.446161e-09, 
    -2.83643e-10, -3.241439e-10, -1.154405e-09, -3.490754e-10, 2.582681e-10, 
    2.685852e-10, 1.503215e-09, 1.181988e-11, -1.602984e-10, 1.250044e-08, 
    -1.962519e-10, 6.330083e-10, 9.795826e-10, 1.145168e-09, -4.850165e-10, 
    -1.608925e-09, 2.088143e-10, -1.236401e-09, -7.547953e-10, 1.27153e-09, 
    1.091394e-12, 9.791279e-12, -6.393641e-11, -4.393641e-11, 9.578116e-11,
  4.203976e-09, -6.109325e-09, -5.314767e-09, -2.122441e-09, -2.204949e-09, 
    6.064695e-10, 4.193147e-09, 2.858663e-09, 3.320402e-09, 5.864202e-09, 
    4.062834e-09, 2.957769e-09, 7.255565e-10, 1.592134e-09, -2.090921e-09, 
    -1.210985e-09, -9.718477e-10, 1.621594e-09, -1.110788e-09, -1.922373e-10, 
    -8.440537e-11, 7.3954e-10, 2.65068e-10, -2.417401e-09, 2.512088e-09, 
    -4.473314e-09, -5.809419e-09, -3.948848e-09, -1.390099e-09, 
    -6.043727e-09, 2.981123e-08, 1.455513e-08, -3.371774e-09, 2.099803e-09, 
    -1.605471e-10, 1.269729e-08, 6.183328e-10, -1.870504e-11, 2.921617e-09, 
    -3.466449e-09, 3.000749e-09, -1.49889e-10, 3.209735e-10, 3.481389e-10, 
    3.056904e-09, 5.987957e-10, -1.422784e-09, -1.665313e-09, -3.801503e-10, 
    -1.685851e-10, 4.637855e-10, -3.594423e-10, 9.296726e-10, -1.175337e-10, 
    -6.11788e-10, -1.175948e-11, -3.579736e-09, 5.440346e-09, -5.808782e-09, 
    6.427214e-10, -7.070611e-11, -2.148894e-10, -5.918466e-10, -7.059482e-10, 
    4.618102e-11, -7.149247e-09, 2.729344e-09, -3.176829e-09, 5.251486e-09, 
    -4.63293e-09, 7.087024e-10, -2.75039e-09, -1.264361e-09, 4.670319e-09, 
    4.279052e-09, -2.084661e-10, 3.26601e-11, 2.990035e-10, 5.228529e-11, 
    2.829502e-09, -1.014378e-09, -4.984201e-10, 4.502709e-11, -2.804574e-08, 
    2.267235e-09, 7.282566e-10, 2.208573e-09, 1.427694e-10, 8.487704e-10, 
    1.821334e-10, -9.026095e-10, 1.818963e-09, 9.733014e-11, 8.505951e-09, 
    -1.732296e-09, -2.525198e-10, -3.864883e-10, -3.937188e-10, -5.22725e-10, 
    4.07654e-10, 5.005134e-10, 1.440068e-09, -1.007194e-12, -2.934843e-10, 
    7.755666e-09, -1.371113e-09, -6.785683e-12, -4.026148e-10, -9.669279e-10, 
    -1.130381e-09, 8.426539e-10, 1.329376e-09, -9.090613e-10, -1.913563e-10, 
    2.017835e-09, -9.619328e-12, 4.461498e-11, -5.683276e-11, -4.446399e-11, 
    4.087752e-11,
  5.365081e-09, -4.914199e-09, -4.560803e-09, -1.555293e-09, -1.788379e-09, 
    -1.719314e-09, 4.335135e-09, 1.474859e-09, 2.259412e-09, 7.614545e-09, 
    1.062162e-08, 6.371124e-09, 1.591559e-09, 5.770062e-09, -2.549996e-09, 
    -2.978509e-10, -1.457033e-09, 1.549637e-09, -1.618549e-09, -9.867449e-10, 
    -7.77618e-11, 7.638334e-10, 4.457092e-10, -2.330921e-09, 1.238311e-08, 
    1.045606e-08, -6.336194e-09, 2.108521e-09, -6.837865e-09, -8.252613e-09, 
    2.587112e-08, 1.391555e-08, 4.427591e-09, 3.804359e-09, -8.412826e-11, 
    1.944349e-08, 1.268373e-09, -2.693454e-10, 8.08808e-09, -2.002537e-09, 
    2.678826e-09, -3.596767e-10, -1.000302e-09, -8.101608e-11, 6.730261e-11, 
    -7.279084e-10, 2.959538e-09, -1.500453e-10, -5.997947e-10, -5.863754e-11, 
    3.836398e-10, -2.029822e-09, 1.752406e-09, -1.199851e-10, -9.22553e-10, 
    -2.259526e-11, -5.057501e-09, 2.907876e-09, -9.554411e-10, 2.03087e-09, 
    -4.795879e-10, -2.54488e-10, -1.40264e-09, 1.036216e-09, -2.7988e-10, 
    -1.107446e-08, 2.855245e-10, -1.718405e-09, 1.16606e-08, -7.452371e-09, 
    3.620926e-10, -2.087319e-09, -1.0414e-09, 4.944496e-09, -6.868193e-10, 
    -1.171259e-10, 5.0278e-11, 4.953833e-10, -2.651106e-11, 4.346504e-09, 
    -1.07724e-09, -3.990792e-10, 9.065531e-10, -2.247788e-09, 1.377231e-09, 
    5.857714e-10, 2.527145e-09, 1.499529e-10, 2.658105e-10, -1.374261e-09, 
    -2.88415e-09, 1.113971e-09, 1.202949e-10, 2.864284e-08, 2.239858e-09, 
    -2.722743e-10, -4.052026e-10, 1.695412e-09, -7.544827e-10, 6.688424e-10, 
    -3.100808e-11, 1.338414e-09, -2.326495e-11, -3.543725e-10, 6.421999e-09, 
    -1.603524e-09, -7.879635e-10, -2.677467e-09, -4.981473e-09, 
    -2.986468e-09, 4.518967e-09, 2.943864e-09, -5.039738e-10, 4.571632e-10, 
    2.86505e-09, -4.646381e-11, 7.97975e-11, 5.047784e-11, -2.35687e-11, 
    -1.009539e-10,
  3.876323e-09, 6.82121e-10, -4.409856e-09, -5.620166e-09, -1.321041e-09, 
    -3.259231e-09, 3.91077e-09, 2.629633e-09, 9.816858e-11, 5.35897e-09, 
    1.342687e-08, 1.080309e-08, -1.534772e-12, -2.722231e-10, 1.421085e-10, 
    1.500156e-10, -1.568787e-09, 7.711947e-10, 1.86003e-09, -2.502304e-09, 
    4.166623e-11, 2.365255e-10, 3.807941e-10, -7.9865e-10, 1.661778e-08, 
    2.605998e-08, -3.491323e-09, 7.406697e-09, -9.833116e-09, -8.682719e-09, 
    2.424463e-08, 1.552604e-08, 9.16566e-09, 4.330502e-09, 1.762146e-11, 
    2.538445e-08, 1.905249e-09, -4.452971e-11, 1.442208e-08, -2.443312e-09, 
    2.784077e-09, -3.188347e-10, -1.659657e-09, -5.975185e-10, 1.191268e-09, 
    -1.860997e-09, 4.312199e-09, -1.670202e-10, -6.905566e-10, 1.08642e-11, 
    7.389218e-10, -2.412094e-09, 2.346962e-09, 5.991296e-12, -1.540866e-09, 
    -6.681944e-11, -6.270056e-09, 4.22192e-09, 6.967693e-10, 2.759442e-09, 
    -8.670327e-10, -5.395577e-10, -2.022716e-09, -6.471625e-10, 
    -5.085212e-10, -3.977846e-09, 3.34569e-09, 2.887134e-09, 2.245565e-08, 
    -1.13381e-08, 9.362111e-11, -1.852641e-09, 9.055157e-10, 8.910774e-10, 
    2.298304e-09, -1.172111e-10, 6.311041e-11, 6.69246e-10, -1.747892e-10, 
    7.852179e-09, -8.770087e-10, 6.498908e-11, 2.352664e-09, 1.55311e-08, 
    2.506795e-09, 1.743956e-09, 1.472813e-09, 2.792717e-10, -4.101359e-10, 
    -4.359606e-09, -6.494929e-09, -1.420641e-10, 5.890399e-11, 3.291974e-08, 
    6.096457e-10, -1.094173e-09, -4.010189e-10, 4.187825e-09, -1.054275e-09, 
    1.017781e-09, -1.198714e-09, 1.043432e-09, -7.930367e-11, -2.812008e-10, 
    8.235475e-10, -7.889298e-10, -7.943299e-10, -4.946457e-09, -6.861683e-09, 
    -3.263153e-09, 1.175619e-08, 3.32426e-09, -4.869776e-10, 1.314959e-09, 
    3.816467e-09, -1.711555e-11, 1.203304e-10, 1.557634e-10, -2.492939e-11, 
    -2.609113e-10,
  2.609795e-09, 1.367823e-09, -6.609753e-10, -8.603251e-10, 4.942535e-10, 
    -3.871151e-09, 2.899014e-09, 5.126992e-09, -8.494681e-10, 3.208243e-09, 
    8.959262e-09, 1.764346e-08, -8.967618e-10, -2.073875e-09, -1.947456e-10, 
    -1.382597e-09, -1.587472e-09, -1.861338e-10, 5.820276e-09, -4.195044e-09, 
    -3.807372e-10, -4.262688e-10, 3.240075e-12, 7.531753e-11, 9.205451e-09, 
    1.747696e-08, -1.595481e-09, 1.210321e-08, 4.331071e-09, -5.92695e-09, 
    2.778279e-08, 1.966487e-08, 1.048898e-08, 4.478864e-09, 4.169465e-10, 
    2.796702e-08, 1.758849e-09, 2.694094e-10, 1.755666e-08, -4.205548e-09, 
    3.91052e-09, -3.175273e-10, -1.789871e-09, -1.373524e-09, 6.217874e-09, 
    2.452794e-09, 9.00809e-09, -7.715641e-10, -9.654059e-10, 3.473133e-11, 
    1.148067e-09, -1.851731e-09, 3.028862e-09, 5.264837e-11, -2.718939e-09, 
    -1.127205e-10, -1.03239e-08, 5.992535e-09, 8.104724e-09, 2.914234e-09, 
    -6.173195e-11, -1.057458e-09, -1.51357e-09, -2.118838e-09, -1.097101e-09, 
    -3.140372e-09, 7.867527e-09, 1.63771e-08, 1.40526e-08, -1.51299e-08, 
    -5.923084e-11, -1.912724e-09, -3.322498e-10, -2.729621e-09, 3.271943e-09, 
    -2.220304e-10, 6.834711e-11, 3.503686e-10, -2.564676e-10, 1.310593e-08, 
    -6.683365e-10, 3.808594e-10, 5.45657e-09, 8.720065e-09, -3.76474e-10, 
    1.389878e-09, 4.240519e-10, 2.320348e-10, -5.331113e-10, -8.231353e-09, 
    -9.061694e-09, -1.738272e-09, -1.307399e-10, 1.366803e-08, -3.964772e-09, 
    -2.963208e-09, -3.596256e-10, 7.962228e-09, -1.339458e-09, 1.412298e-09, 
    1.736225e-09, -6.256329e-10, -2.457838e-10, -1.298908e-10, 8.525433e-09, 
    -1.081162e-10, -2.266916e-10, -2.205013e-09, -4.379331e-09, 2.905097e-09, 
    1.70059e-08, 2.723425e-09, -1.380499e-09, 2.508159e-09, 4.715275e-09, 
    -4.89365e-11, 1.45306e-10, 1.836717e-10, -4.077449e-11, -3.246896e-10,
  1.959961e-09, 1.458091e-09, 1.49771e-09, 1.415344e-09, 1.227363e-09, 
    -3.531511e-09, 1.765045e-09, 5.518871e-09, 1.380556e-09, 2.802153e-09, 
    5.899665e-09, 1.423189e-08, -5.329071e-10, -9.118253e-10, 3.970342e-09, 
    -3.235738e-09, -3.984269e-10, -2.688552e-09, 1.161142e-08, -6.275286e-09, 
    -5.261768e-09, -6.083951e-10, 5.144329e-11, 9.397922e-10, 1.394653e-09, 
    2.870252e-09, -2.652541e-09, 1.638199e-08, 1.1118e-08, 9.820269e-10, 
    2.972916e-08, 2.701523e-08, 1.110425e-08, 7.160054e-09, -9.429755e-10, 
    2.657333e-08, 2.337686e-10, 3.455725e-10, 1.881091e-08, -3.994545e-09, 
    6.352309e-09, -7.257199e-10, -2.242444e-09, -2.045108e-09, 1.970932e-09, 
    4.274511e-09, 9.225829e-09, -5.597798e-10, -2.830552e-09, 7.293721e-11, 
    1.324764e-09, -1.041542e-09, 3.794321e-09, 2.758043e-11, -4.906049e-09, 
    -9.160317e-11, -1.487558e-08, 7.858068e-09, 1.803846e-08, 2.707594e-09, 
    2.674369e-09, -1.639478e-09, -6.515961e-10, -4.150809e-09, -3.173432e-09, 
    -5.726577e-09, 4.566937e-08, 4.158539e-08, 4.250637e-09, -1.468186e-08, 
    6.82121e-13, -3.341142e-09, -5.455263e-09, -8.868142e-10, 9.954825e-09, 
    -2.340244e-10, 7.703704e-11, -1.477503e-10, -3.730193e-10, 1.526615e-08, 
    -1.305409e-09, -3.751296e-10, 1.000799e-08, 2.135039e-09, -4.304013e-09, 
    1.620947e-09, 9.061409e-10, 3.075229e-11, -2.113101e-10, -1.479737e-08, 
    -4.219942e-09, -3.209003e-09, -3.332872e-10, -9.73896e-09, -8.514405e-09, 
    -5.434265e-09, -3.778609e-10, 1.083316e-08, -1.259082e-09, 1.85936e-09, 
    3.074433e-09, -4.325425e-09, -5.724665e-10, -3.968381e-11, 1.673988e-08, 
    -2.142997e-11, 8.578809e-10, -5.214815e-10, -3.554533e-09, 2.986042e-09, 
    1.571783e-08, 7.107133e-10, -3.907701e-09, 4.746653e-09, 4.127855e-09, 
    -4.468461e-11, 1.564402e-10, 2.355947e-10, -5.722356e-11, -1.253397e-10,
  -1.871854e-10, 1.749981e-09, 3.022933e-10, 1.555293e-09, 1.725994e-09, 
    -7.138965e-10, 5.671268e-10, 4.067317e-09, 1.634362e-09, -8.795382e-10, 
    6.468611e-09, 1.401708e-08, 2.16545e-09, 1.566377e-09, 5.938091e-09, 
    -1.765966e-09, 1.938866e-09, -6.35734e-09, 2.007936e-08, -8.429708e-09, 
    -1.423291e-08, -4.702088e-10, 1.186152e-09, 1.275396e-09, -5.792344e-10, 
    5.504717e-10, -7.287326e-11, 1.26397e-08, 1.680786e-08, -1.476792e-09, 
    3.097682e-08, 3.933735e-08, 1.190369e-08, 1.270325e-08, -8.907364e-09, 
    2.769303e-08, 1.458096e-09, 4.820322e-10, 1.579599e-08, -4.093167e-09, 
    8.319955e-09, -2.665388e-10, 9.510899e-10, -2.368897e-09, -6.241407e-09, 
    2.970739e-08, 6.804981e-09, 2.506511e-10, -8.13917e-09, 1.437535e-10, 
    -5.578187e-10, 2.016236e-09, 3.948145e-09, -1.350713e-10, -7.455263e-09, 
    -5.115908e-13, -1.434591e-08, 1.412497e-08, 6.11301e-09, 1.745285e-09, 
    3.386674e-09, -3.232458e-09, 2.506226e-10, -4.604135e-09, -7.077256e-09, 
    4.254844e-09, 9.304222e-08, 6.308545e-08, 2.658055e-09, -6.814787e-09, 
    4.800995e-10, 2.648903e-09, -3.877176e-09, 8.855068e-10, 1.484615e-08, 
    -2.38515e-10, 1.927063e-10, 3.680469e-10, -3.760604e-10, 1.71496e-08, 
    -4.189133e-09, -1.702018e-09, 1.565189e-08, 3.000991e-09, -3.466653e-09, 
    -2.383956e-09, 4.112735e-09, -4.071126e-10, 3.449935e-09, -2.404727e-08, 
    8.847962e-09, -4.080711e-09, -7.753442e-11, -1.179507e-08, -8.345694e-09, 
    -6.808739e-09, -4.905473e-10, 8.550558e-09, -3.270202e-10, 2.501895e-09, 
    1.938474e-09, -6.279432e-09, -6.06093e-10, -1.795186e-11, 1.926242e-08, 
    -4.174922e-09, 2.433467e-09, 4.855565e-10, -7.603376e-10, 7.267886e-09, 
    1.15233e-08, 9.29731e-10, -7.095025e-09, 9.572602e-09, 3.916341e-09, 
    -2.80238e-12, 1.385558e-10, 3.544489e-10, -7.235457e-11, -1.311946e-10,
  3.531682e-10, 2.270497e-09, -4.371827e-10, -1.351737e-10, 1.819444e-09, 
    4.534968e-10, -1.376634e-09, 4.248932e-09, -9.379164e-11, -1.490548e-09, 
    9.524683e-10, 1.132616e-08, 1.325759e-09, 1.631332e-08, -3.492289e-09, 
    -1.337713e-09, 4.250813e-09, -1.468882e-08, 2.685299e-08, -5.015977e-09, 
    -1.684776e-08, -1.032788e-09, 3.006619e-09, 9.055157e-11, -4.662866e-10, 
    2.950742e-10, 1.373718e-08, -1.12891e-09, 1.726119e-08, 2.862635e-09, 
    3.273522e-08, 5.432025e-08, 1.331006e-08, 1.525177e-08, -1.908592e-08, 
    3.536371e-08, -3.726882e-10, 4.418084e-10, 5.401546e-09, -5.555997e-09, 
    7.41353e-09, 2.680622e-09, 8.120523e-09, -2.276924e-09, -5.411323e-09, 
    4.318889e-08, 1.208466e-08, 1.739636e-09, -1.661781e-08, 2.135891e-10, 
    -3.3668e-09, 3.244622e-10, 7.144275e-09, -3.644118e-10, -6.936972e-09, 
    1.798526e-10, -1.48425e-08, 2.463588e-08, -2.706078e-08, 2.812591e-09, 
    8.217285e-10, -9.055498e-09, 7.418635e-10, -4.671972e-09, -1.116465e-08, 
    6.909204e-09, 6.49855e-08, 6.544167e-08, -1.004537e-09, 8.402594e-10, 
    1.017497e-10, 1.234929e-08, 3.114508e-09, 7.067911e-10, 1.848328e-08, 
    -2.015668e-10, 2.84416e-10, -1.53193e-10, 2.663536e-11, 2.00032e-09, 
    -8.672174e-09, -8.328925e-10, 2.319427e-08, 1.094804e-09, 6.671769e-09, 
    -4.771834e-09, 9.209771e-10, 1.447802e-09, 4.265969e-09, -2.815767e-08, 
    1.081082e-08, -3.726747e-09, -2.90953e-10, 3.826051e-09, -8.428856e-09, 
    -7.648339e-09, -8.33586e-10, -2.133504e-09, 1.837805e-09, 3.464606e-09, 
    -3.731202e-10, 5.976233e-10, -9.196555e-11, -2.771223e-10, 1.354363e-08, 
    5.137281e-09, 5.595382e-09, -4.362846e-09, 1.665285e-09, 5.005006e-09, 
    6.014432e-09, -2.516458e-10, -4.32658e-09, 1.367829e-08, 5.208619e-09, 
    -8.290044e-11, 5.988454e-11, 5.047855e-10, -5.405809e-11, -7.960352e-10,
  -2.441425e-10, 7.243557e-10, 3.745868e-09, 8.823804e-10, 2.652143e-09, 
    5.189804e-11, -7.78283e-09, 6.682285e-09, -1.240778e-09, 1.300236e-09, 
    -2.905495e-09, 7.7506e-10, -2.43989e-09, 4.210068e-08, -3.363084e-09, 
    -5.838922e-09, 6.112015e-09, -2.243686e-08, 2.771083e-08, 2.074898e-09, 
    -1.071413e-08, -1.109811e-09, 4.116089e-09, -1.917897e-09, 2.012825e-09, 
    2.59638e-09, 2.047216e-08, -1.455902e-08, -1.76334e-09, 8.203813e-09, 
    3.805701e-08, 7.259689e-08, 1.32614e-08, 1.774066e-08, -1.857762e-08, 
    4.158989e-08, 8.894063e-10, 9.130474e-10, -1.003241e-08, -7.220308e-09, 
    3.190053e-09, 5.532002e-10, 1.193001e-08, -1.534561e-09, -1.566968e-08, 
    3.701831e-08, 2.172672e-08, 2.298492e-09, -2.641939e-08, 3.248033e-10, 
    -6.843919e-09, -2.44853e-09, 1.328513e-08, -7.981612e-10, -2.427691e-09, 
    4.525873e-10, -2.049222e-08, 3.617129e-08, -3.526212e-08, -3.97668e-09, 
    -8.859047e-09, -1.475178e-08, 4.626486e-10, -7.179755e-09, -1.534017e-08, 
    1.221144e-08, 6.627027e-08, 6.192255e-08, 8.339327e-09, 3.372577e-09, 
    -2.030276e-09, 2.250545e-09, -1.336304e-08, 5.295192e-09, 2.390144e-08, 
    -9.691803e-11, 4.64091e-10, -5.502727e-10, 2.537909e-09, -1.149374e-09, 
    -1.15779e-08, -2.858773e-09, 2.925592e-08, 1.986109e-10, 6.451842e-09, 
    -3.419927e-09, -1.189511e-08, -3.597052e-10, 5.14234e-09, -3.00021e-08, 
    2.006345e-09, 1.929585e-10, -2.845979e-09, 5.685344e-09, -1.310167e-08, 
    -7.121281e-09, -3.094328e-10, -1.493822e-08, 4.932303e-09, 4.504693e-09, 
    1.203944e-10, 1.107533e-08, 7.604619e-10, -1.079222e-09, 1.889924e-08, 
    6.723099e-09, 1.754586e-09, -7.781068e-09, -1.222134e-11, 2.122249e-09, 
    2.818524e-09, -3.60933e-09, 5.199468e-10, 1.794757e-08, 4.346418e-09, 
    -2.174204e-10, -1.996625e-11, 6.138272e-10, -4.749623e-11, -8.517418e-10,
  -4.471872e-10, -2.131401e-09, 2.055936e-08, 6.124935e-09, 5.112724e-09, 
    -1.915112e-09, -1.420381e-08, 5.777622e-09, 2.005265e-09, 2.178297e-09, 
    2.160618e-10, -1.798298e-09, 1.58866e-09, 8.670611e-09, 3.074706e-08, 
    -1.436438e-08, 6.916145e-09, -3.221578e-08, 2.521778e-08, 6.589403e-09, 
    -2.576428e-09, -2.74639e-09, 3.050104e-09, -2.869569e-09, 4.148148e-09, 
    3.140144e-09, 5.083308e-08, -1.818091e-08, -6.067512e-08, 2.177484e-08, 
    4.743339e-08, 8.709355e-08, 1.370842e-08, 2.856586e-08, -7.080132e-09, 
    4.338807e-08, -1.048448e-09, 1.567734e-09, -3.138075e-08, -1.67346e-08, 
    -3.147909e-09, -1.545573e-09, 1.302487e-08, -7.824212e-10, -2.075723e-08, 
    1.237424e-08, 2.519269e-08, -4.369795e-09, -3.169805e-08, 4.684928e-10, 
    -1.231328e-08, -3.153559e-09, 1.595721e-08, -2.070203e-09, -3.142337e-09, 
    6.009486e-10, -4.379496e-08, 4.954353e-08, -4.901477e-09, -1.965506e-08, 
    -1.100932e-08, -1.663182e-09, -8.237748e-10, -8.663721e-09, 
    -2.018412e-08, 2.645589e-08, 2.4531e-08, 5.959811e-08, 5.240224e-09, 
    1.615263e-09, -2.035222e-09, -1.921438e-08, -5.373937e-08, 9.638654e-09, 
    3.175518e-08, 1.966214e-10, 9.42677e-10, -1.736112e-09, 8.555236e-09, 
    3.59783e-08, -1.872004e-08, -3.079086e-08, 2.755647e-08, 2.399929e-09, 
    -1.334968e-09, 8.323013e-10, -1.906847e-08, -8.498034e-09, 2.619873e-09, 
    -3.409625e-08, 1.182343e-10, 7.575661e-09, -6.379196e-09, 6.114931e-11, 
    -1.906011e-08, -2.846497e-09, 7.906943e-09, -1.604661e-08, 6.034441e-09, 
    4.885442e-09, 7.47832e-10, 1.55153e-08, 1.57592e-09, -1.35152e-09, 
    2.393762e-08, -1.072863e-09, -4.03827e-09, -8.365078e-10, 1.178478e-09, 
    1.294154e-09, 1.645731e-09, -5.678146e-09, 2.728541e-09, 1.753392e-08, 
    -2.951879e-10, -4.111484e-10, 8.875389e-11, 6.57792e-10, -2.648548e-11, 
    -1.627598e-09,
  -2.726097e-09, 1.028297e-10, 4.046683e-08, -4.073399e-10, 7.695405e-09, 
    -2.398679e-09, -1.194275e-08, 1.488218e-09, 4.179185e-09, 3.373771e-09, 
    2.537092e-09, -2.105594e-09, 1.241574e-09, 8.429879e-11, 1.594634e-08, 
    -2.721814e-08, 7.52641e-09, -4.405243e-08, 2.335077e-08, 1.120799e-08, 
    8.154188e-10, -1.221792e-08, -1.668639e-09, -2.147772e-09, 3.434138e-09, 
    2.13771e-09, 8.540525e-08, -1.954027e-08, -8.672475e-08, 3.499713e-08, 
    4.866524e-08, 9.600791e-08, 1.141348e-08, 4.649195e-08, -2.058755e-09, 
    5.101759e-08, -1.849889e-09, 1.979942e-09, -5.908259e-08, -3.381958e-08, 
    -1.797157e-08, 1.013973e-09, 1.415903e-08, -1.1604e-09, -2.127717e-08, 
    6.141534e-09, 3.432078e-08, -1.982724e-08, -2.705934e-08, 5.209593e-10, 
    -1.946774e-08, -4.073058e-09, 1.332036e-08, -2.249647e-09, -1.563158e-08, 
    6.569394e-10, -7.737447e-08, 6.423958e-08, 5.466191e-08, -1.932052e-08, 
    -1.340641e-08, 4.847493e-09, 9.742962e-11, -1.106996e-08, -2.39715e-08, 
    1.527576e-08, -1.620037e-09, 5.822181e-08, 1.469664e-08, 1.380658e-08, 
    -1.997876e-09, -3.078191e-08, -6.466485e-08, 4.479205e-09, 3.819784e-08, 
    7.70342e-10, 9.226113e-10, -3.596384e-09, 1.222188e-08, 5.271062e-08, 
    -2.411582e-08, -8.922309e-08, 1.859308e-08, 2.207514e-09, -6.559731e-10, 
    2.701427e-09, -9.611313e-09, -1.191148e-08, 2.544407e-09, -4.010349e-08, 
    2.540901e-11, 1.615039e-08, -6.276238e-09, 1.078035e-08, -2.197362e-08, 
    -7.236395e-09, 3.048704e-08, 2.943636e-09, 4.024741e-09, 3.891864e-09, 
    -1.425633e-10, 8.879439e-09, -1.523279e-09, -1.340091e-09, 2.256076e-08, 
    -8.946813e-09, -2.209731e-09, 7.717347e-09, 4.181118e-09, 1.446097e-09, 
    4.117737e-10, -9.96522e-10, 2.973536e-09, 1.047397e-08, -9.969256e-09, 
    -6.446612e-10, 7.363354e-10, 9.169181e-10, -3.975487e-12, -5.047696e-09,
  4.738035e-08, 3.653895e-09, 5.377194e-08, -1.277976e-08, 1.077342e-08, 
    -1.44837e-09, -4.944013e-09, -2.221782e-09, 2.842057e-09, 5.596348e-09, 
    1.754984e-09, 3.611831e-10, 6.82121e-13, -3.581818e-09, -5.884999e-09, 
    -3.735208e-08, 7.685446e-09, -5.905412e-08, 1.903568e-08, 2.797685e-08, 
    -6.899086e-09, -2.053332e-08, -2.755201e-09, -1.567059e-09, 1.678814e-09, 
    1.14278e-09, 1.323241e-07, -1.669457e-08, -2.953425e-08, 4.270828e-08, 
    4.649155e-08, 7.549727e-08, -6.057235e-10, 5.78076e-08, -1.162618e-08, 
    7.68465e-08, -1.770741e-09, 2.870834e-09, -8.15777e-08, -4.755157e-08, 
    -3.186528e-08, 3.31886e-09, 1.282996e-08, -1.846276e-09, -9.120754e-09, 
    3.496621e-08, 3.95828e-08, -2.764938e-08, -2.616891e-08, 4.205916e-10, 
    -2.509906e-08, -7.663516e-09, 2.211398e-08, -3.738524e-09, -2.576841e-08, 
    4.45425e-10, -9.925122e-08, 7.609221e-08, 1.181828e-07, -2.798367e-08, 
    -1.186686e-08, 5.474476e-09, 4.171284e-09, -1.11173e-08, -2.688212e-08, 
    4.320418e-08, 4.867729e-09, 4.529693e-08, 2.273691e-08, 4.891763e-08, 
    8.966367e-09, -4.185927e-08, -6.375421e-08, -4.180038e-09, 4.306635e-08, 
    1.435524e-09, -1.062674e-09, -6.934357e-09, 1.380706e-08, 3.333741e-08, 
    -2.768672e-08, -1.035416e-07, 1.081673e-08, 2.166871e-09, -6.221171e-09, 
    6.763003e-09, -5.285301e-09, -3.535774e-09, 3.279997e-09, -3.767752e-08, 
    -1.164267e-09, 2.011209e-08, -2.950628e-09, 5.160528e-08, -2.147851e-08, 
    -2.199134e-08, 6.167101e-09, 9.616429e-09, 1.195644e-09, 1.708349e-09, 
    -1.945182e-10, 2.013202e-09, -6.762086e-09, -1.953488e-09, 3.89025e-08, 
    -1.238686e-08, -4.949811e-09, 4.764047e-09, 7.219796e-09, 5.968559e-10, 
    1.523517e-09, 5.762786e-10, 7.729568e-10, 4.431058e-09, -2.078082e-08, 
    -8.40123e-10, 1.548301e-09, 8.938343e-10, 3.850431e-11, -6.217988e-09,
  1.792881e-07, 3.676746e-09, 7.090034e-08, -6.844061e-09, 1.650062e-08, 
    -4.428102e-10, 9.097221e-10, -7.626909e-09, 2.44188e-09, 3.260425e-09, 
    1.664375e-09, 2.91675e-09, -1.019089e-09, -1.682474e-08, 9.757741e-10, 
    -4.134627e-08, 7.034146e-09, -5.584184e-08, 1.418583e-08, 4.637195e-08, 
    -1.071658e-08, -7.112931e-09, -7.906124e-09, 1.139711e-09, 4.373533e-10, 
    -8.743655e-10, 1.734895e-08, 4.102048e-09, -1.46282e-08, 4.752155e-08, 
    1.979481e-08, 2.95405e-08, 6.986056e-09, 3.900516e-08, -1.829733e-08, 
    9.984967e-08, -2.534296e-09, 1.707733e-09, -8.082679e-08, -5.516844e-08, 
    -3.255482e-08, 5.668994e-09, 9.662585e-09, -2.99643e-09, 3.329774e-09, 
    4.869821e-08, 4.829019e-08, -3.634335e-08, -1.974411e-08, 1.631832e-10, 
    -2.881922e-08, -2.554452e-08, 1.652482e-08, -5.427591e-09, -2.040585e-08, 
    -1.072635e-10, -9.38079e-08, 8.20768e-08, 2.070624e-07, -5.024491e-08, 
    6.286882e-09, 6.615664e-09, 5.725838e-09, -1.35738e-08, -3.06216e-08, 
    9.712539e-08, -2.93079e-08, 1.687863e-08, 1.736623e-08, 6.307732e-08, 
    3.470961e-08, -6.006144e-08, -4.434378e-08, -5.237325e-09, 4.081861e-08, 
    1.719627e-09, -1.566008e-09, -1.340462e-08, 1.511619e-08, 2.928346e-09, 
    -3.964254e-08, -7.215593e-08, 6.942116e-09, 7.756853e-10, -1.23008e-08, 
    1.462695e-09, 2.866159e-09, 4.834646e-09, 4.953833e-10, -2.767206e-08, 
    -1.007948e-09, 1.37259e-08, -4.154685e-10, 1.599934e-07, -1.484545e-08, 
    -1.66737e-08, -2.121744e-08, 1.290709e-08, -2.72621e-09, -7.206836e-10, 
    6.830305e-10, 7.475833e-10, -2.400917e-09, -1.504063e-09, 9.108999e-08, 
    -1.364924e-08, -1.311105e-08, 1.930403e-09, 1.081139e-08, -4.813501e-10, 
    1.364697e-09, 1.204626e-09, -1.617764e-10, -5.976517e-10, -1.570913e-08, 
    -1.16695e-09, 2.63698e-09, 5.679581e-10, 2.426503e-11, -2.713591e-09,
  1.388614e-07, 1.508681e-09, 8.66068e-08, -8.020436e-09, 2.355188e-08, 
    3.929756e-09, -5.969127e-10, -7.950746e-09, -3.326079e-09, 1.966214e-10, 
    1.6949e-09, 3.123603e-09, 8.918732e-11, -3.33153e-08, 3.18704e-09, 
    -4.553689e-08, 4.208084e-09, -4.736052e-08, 1.616378e-08, 3.753729e-08, 
    -1.12189e-08, 3.606431e-09, -1.947507e-08, 6.317066e-09, 2.385889e-09, 
    -7.33138e-09, -4.061343e-08, 1.931937e-09, -2.933388e-08, 2.956045e-08, 
    -8.096151e-09, -3.448071e-08, 2.435746e-08, 2.844234e-08, -1.688562e-08, 
    9.116189e-08, -1.463081e-09, -2.268507e-09, -1.189636e-08, -6.094594e-08, 
    -2.229739e-08, 9.047938e-09, 1.115743e-08, -6.056233e-09, 5.860386e-09, 
    4.238217e-08, 6.581172e-08, -5.65808e-08, -5.103641e-09, -3.04496e-10, 
    -3.211861e-08, -4.823829e-08, -1.504463e-08, -7.163828e-09, 
    -1.034181e-08, -5.537117e-10, -7.688328e-08, 9.614534e-08, 2.884104e-07, 
    -7.375468e-08, 1.02844e-08, 4.248761e-09, 7.302049e-09, -1.709544e-08, 
    -2.75351e-08, 6.896909e-08, -5.710268e-08, 5.835716e-09, 1.694156e-08, 
    -8.466202e-09, 2.476889e-08, -7.038324e-08, -5.590147e-08, 9.602559e-10, 
    3.002599e-08, 1.257888e-09, -1.930928e-09, -2.398147e-08, 1.566694e-08, 
    -5.049452e-08, -4.43053e-08, -5.300859e-08, 4.629499e-09, -5.912113e-09, 
    -2.712625e-09, -5.920691e-08, 1.534369e-08, 3.339153e-09, 8.965145e-09, 
    -2.398002e-08, -2.336265e-11, 3.803223e-09, -3.525997e-10, 2.615036e-07, 
    -2.106248e-08, 2.156991e-08, -1.064005e-08, 1.607253e-08, -5.339587e-09, 
    -3.287903e-09, 4.278661e-09, -4.675655e-10, 4.940823e-09, 2.283258e-10, 
    4.017335e-08, -2.658061e-08, -2.088512e-08, -2.787033e-10, 1.376367e-08, 
    -3.639684e-10, -4.231993e-10, 1.020169e-09, -5.999823e-10, -1.733213e-09, 
    -1.421597e-09, -2.595527e-09, 3.367333e-09, 3.330349e-10, -3.746692e-11, 
    5.071058e-09,
  2.323657e-08, 2.437446e-10, 8.16417e-08, -6.391713e-08, 2.322747e-08, 
    1.904834e-08, -3.265427e-09, -3.750529e-09, -6.348841e-09, 3.133437e-09, 
    4.095909e-09, 2.083084e-09, -1.801368e-09, -4.898584e-08, 7.706035e-09, 
    -4.699577e-08, -4.314757e-09, -3.946712e-08, 2.308124e-08, 1.064291e-08, 
    -1.65345e-08, 7.094059e-10, -2.477691e-09, 1.15341e-08, -4.874551e-09, 
    -6.022333e-09, -1.035165e-07, -1.774879e-08, -1.901572e-08, 1.390379e-08, 
    -1.087687e-08, -7.337667e-08, 2.352715e-08, 3.109881e-08, -1.580554e-08, 
    6.133405e-08, 1.470084e-10, -5.001212e-09, 4.169351e-09, -6.692404e-08, 
    -1.18107e-08, 8.879397e-09, 1.172833e-08, -5.905916e-09, 1.484523e-09, 
    4.435742e-08, 6.533469e-08, -3.763961e-08, 5.518313e-09, -1.344283e-09, 
    -3.181765e-08, -6.662117e-08, -4.667357e-08, -1.055141e-08, 
    -5.078101e-09, -1.369926e-10, -6.321409e-08, 1.21136e-07, 3.193409e-07, 
    -8.848824e-08, 2.434945e-09, 2.460638e-09, 3.584319e-09, -3.012208e-08, 
    -1.125932e-08, 6.619905e-08, 7.387371e-10, 1.42586e-08, 1.300157e-08, 
    -6.05587e-09, 4.749666e-08, -9.365635e-08, -7.557242e-08, 1.086403e-08, 
    2.526876e-08, -2.363549e-10, -2.544581e-09, -3.89627e-08, 1.540533e-08, 
    -5.3848e-08, -5.206294e-08, -5.537972e-08, 4.011042e-09, -9.337555e-09, 
    7.522431e-09, -9.703774e-08, 8.284246e-09, 1.100375e-09, 1.566533e-08, 
    -2.396018e-08, -1.684271e-09, 7.685941e-10, -1.690097e-09, 3.375289e-07, 
    -3.259299e-08, 6.222035e-08, -5.489369e-09, 2.403056e-08, -5.420702e-09, 
    -7.128961e-09, 3.444507e-08, -1.105858e-08, 1.3425e-08, 1.757392e-09, 
    -5.619506e-08, -1.932756e-08, -2.804268e-08, -3.917648e-10, 1.938952e-08, 
    1.685976e-10, -2.04227e-09, 9.049472e-11, -2.288971e-09, -1.230546e-09, 
    1.218609e-09, -3.380558e-09, 3.129372e-09, 3.594174e-10, -1.160245e-10, 
    -2.814886e-10,
  -4.781157e-08, -3.080913e-11, 4.44021e-08, -8.981624e-08, 4.057392e-08, 
    2.614809e-08, -9.106316e-09, 8.396114e-09, -7.323706e-09, 4.558842e-09, 
    8.446932e-10, -9.430323e-10, -4.321691e-09, -8.421694e-08, 9.206474e-09, 
    -4.428331e-08, -8.116182e-09, -3.613673e-08, 2.508784e-08, -2.787715e-09, 
    -1.85272e-08, 3.520313e-08, 1.244985e-09, -2.848424e-09, -6.37101e-09, 
    2.082743e-09, -5.244863e-08, -2.810884e-08, -2.155275e-09, 1.071498e-08, 
    3.61149e-09, -5.970651e-08, 4.954813e-09, -1.912167e-08, -1.91568e-08, 
    3.6443e-08, 1.438548e-09, -6.165635e-09, -2.181082e-09, -6.424932e-08, 
    -2.410263e-08, 5.550874e-09, 3.914977e-09, -1.641045e-09, -6.206392e-09, 
    3.949458e-08, 7.043241e-08, -1.642394e-08, 7.480185e-09, -1.894257e-09, 
    -2.956851e-08, -5.980553e-08, -7.650328e-08, -1.171954e-08, 1.312667e-09, 
    1.961098e-10, -7.193046e-08, 1.483092e-07, 2.981161e-07, -6.730082e-08, 
    6.306209e-10, 8.889174e-10, 1.5909e-08, -6.425716e-08, 9.836413e-09, 
    5.046127e-08, 2.544016e-08, 2.411821e-08, 1.014246e-08, 2.334093e-08, 
    1.411615e-08, -8.124471e-08, -4.960862e-08, 9.350856e-09, 5.325104e-08, 
    -1.974627e-09, -2.062649e-09, -5.447814e-08, 1.561369e-08, -5.116021e-08, 
    -6.987892e-08, -7.317068e-08, 4.28355e-09, -6.193773e-09, 4.01883e-10, 
    -6.553023e-08, 1.599244e-08, -2.44313e-10, 1.95639e-08, -2.700847e-08, 
    -3.824198e-09, 2.372958e-08, -3.046239e-09, 3.440294e-07, -3.512457e-08, 
    7.006721e-08, -8.900861e-09, 6.089886e-08, -3.406171e-09, -1.218878e-08, 
    2.558875e-08, -1.320637e-08, 1.387264e-08, 5.526957e-10, -6.337348e-08, 
    -1.122226e-08, -3.531272e-08, 1.76658e-09, 3.184755e-08, 9.359269e-09, 
    -1.914714e-09, 7.75799e-10, -2.94051e-09, -1.275907e-09, -1.694275e-09, 
    -4.580522e-09, 3.16561e-09, 3.926104e-11, -1.994849e-10, -1.025307e-08,
  -2.784475e-08, -3.601599e-10, 9.27912e-09, -3.799846e-08, 5.219408e-08, 
    2.209913e-08, -6.283585e-09, 1.025739e-08, 7.449785e-09, 2.910383e-11, 
    1.076614e-10, -7.64885e-10, 5.184575e-09, -8.716847e-08, -1.388582e-08, 
    -3.845706e-08, -2.218153e-08, -3.04014e-08, 1.868189e-08, 3.182208e-09, 
    -2.187915e-08, 9.46718e-08, 1.215494e-08, -1.495812e-08, 2.888214e-09, 
    5.658876e-09, -2.506715e-08, -2.477645e-08, 9.094947e-13, 1.026422e-08, 
    -3.358878e-09, -3.893638e-08, -7.756853e-09, -3.619766e-08, 
    -2.743593e-08, 1.115211e-08, 1.092678e-09, -7.175345e-09, -1.370552e-08, 
    -3.284654e-08, 1.249491e-08, 4.034746e-09, -7.148628e-10, -1.242627e-09, 
    -1.005003e-08, 1.347109e-08, 1.258716e-07, 2.474508e-08, 6.639925e-09, 
    -1.948329e-09, -2.989049e-08, -5.053971e-08, -6.213812e-08, 
    -1.354704e-08, 1.49571e-08, -4.433787e-11, -1.018111e-07, 1.677426e-07, 
    2.026278e-07, -3.561055e-08, -6.82121e-13, 1.47736e-09, 2.009403e-08, 
    -1.013426e-07, 1.03867e-08, 5.372203e-08, 3.815899e-08, 2.756462e-08, 
    3.840682e-09, 2.977094e-08, -2.280084e-07, 1.279886e-09, -3.847799e-08, 
    5.193101e-09, 9.979631e-08, -1.504645e-09, -7.356675e-10, -6.632871e-08, 
    1.690971e-08, -5.600202e-08, -6.348949e-08, -8.321081e-08, 3.43465e-09, 
    -1.253738e-09, -7.066774e-10, -4.732078e-08, -2.938577e-09, 
    -2.073079e-09, 2.343108e-08, -3.110068e-08, 1.774868e-08, 8.483637e-08, 
    -4.048871e-09, 3.194535e-07, -2.213324e-08, 4.430171e-08, -2.063843e-08, 
    5.150468e-08, -6.728214e-09, -2.299637e-08, -2.50958e-08, 5.596661e-10, 
    5.673208e-09, -1.959961e-09, -3.030686e-08, -3.410378e-09, -3.136267e-08, 
    1.22875e-08, 3.190371e-08, 2.230786e-08, -1.206899e-09, -9.068799e-10, 
    -1.965986e-09, -2.85263e-09, -1.884473e-09, -6.025163e-09, 1.814996e-09, 
    -2.08118e-10, -2.924452e-10, 7.877361e-10,
  4.243986e-09, -8.487291e-10, 3.046296e-09, 1.259065e-08, 4.570478e-08, 
    1.946563e-08, -4.017068e-09, 9.643998e-09, 1.540849e-08, 5.883294e-11, 
    -4.543494e-10, 2.051991e-09, 1.847587e-08, -1.862776e-08, 5.65268e-09, 
    -3.096249e-08, -3.942722e-08, -1.143388e-08, -6.005877e-09, 8.500194e-09, 
    3.646505e-10, 1.330783e-07, 7.248713e-08, 9.545317e-09, 7.519304e-09, 
    9.093242e-10, -3.092799e-08, -1.890265e-08, 7.742358e-09, 2.962054e-09, 
    -2.374355e-08, -3.527435e-08, -7.127426e-09, 9.943562e-09, -3.831093e-08, 
    -1.263589e-08, 3.660978e-09, -5.937494e-09, -1.206166e-08, -6.756704e-09, 
    2.87098e-08, 6.191669e-09, -2.414254e-09, -3.871888e-09, 8.571021e-09, 
    -1.428003e-08, 1.479334e-07, 5.554139e-08, 9.465509e-09, -1.321624e-09, 
    -2.849735e-08, -4.355223e-08, 1.633426e-08, -1.625623e-08, 2.937912e-08, 
    -1.003684e-09, -1.284583e-07, 1.957056e-07, 1.047318e-07, -1.704115e-08, 
    9.871997e-10, -9.591247e-09, -1.843563e-08, -1.046233e-07, -3.511706e-08, 
    6.81884e-08, 2.484904e-08, 2.333928e-08, -5.417235e-09, 4.249063e-08, 
    -2.052287e-07, 8.419948e-08, -6.967144e-08, 1.090274e-08, 1.530616e-07, 
    2.029878e-10, 1.679211e-09, -6.593211e-08, 2.017136e-08, -9.880495e-08, 
    -5.280413e-08, -8.118255e-08, -5.676156e-09, -1.64448e-10, -4.16145e-09, 
    -2.915448e-08, -6.048543e-08, -3.907019e-09, 2.595215e-08, -1.115665e-07, 
    8.312435e-08, 1.838892e-07, -6.114476e-09, 2.922602e-07, -6.15313e-09, 
    1.883556e-08, -3.026959e-08, 2.573017e-09, -1.007646e-08, -3.643328e-08, 
    -1.245961e-07, 9.888232e-09, 2.977409e-09, -8.733586e-09, -2.506118e-08, 
    1.968448e-08, -1.077916e-08, 9.383086e-09, 1.740381e-08, 3.538997e-08, 
    9.394512e-10, -3.477055e-09, -3.583693e-09, -5.526715e-09, -1.779824e-09, 
    -6.463688e-09, -2.387281e-09, -2.11184e-10, -3.977334e-10, -1.822156e-08,
  1.379948e-08, -1.763681e-09, 4.243759e-09, 3.057772e-08, 2.3925e-08, 
    2.293865e-08, 1.045549e-08, 9.935718e-09, 1.489587e-08, 5.749087e-09, 
    -3.001844e-09, 1.08156e-09, 2.17654e-08, 5.132034e-08, -7.369692e-09, 
    -2.023523e-08, -4.253286e-08, 2.930403e-08, -1.117803e-07, 9.326243e-09, 
    3.161193e-08, 4.078719e-07, 1.23832e-07, 1.952338e-08, 1.182173e-09, 
    -1.003229e-09, -4.043653e-08, -2.468738e-08, 2.955568e-08, -2.776125e-08, 
    -4.343048e-08, -3.108818e-08, -3.545608e-09, -2.661289e-08, 
    -5.605187e-08, 9.714256e-09, -2.653303e-09, -4.982468e-09, -2.179155e-08, 
    -2.321403e-08, -1.558566e-08, 5.708728e-09, -4.896322e-09, -6.895746e-09, 
    4.218572e-08, -3.275528e-08, 1.211502e-07, 1.101913e-07, 1.827719e-08, 
    -7.399876e-10, -2.305069e-08, -3.108556e-08, 1.028945e-07, -1.804364e-08, 
    4.745505e-08, -2.855245e-09, -1.330854e-07, 2.327022e-07, 8.211818e-08, 
    -8.329209e-09, 2.40351e-09, -5.949704e-08, -1.726579e-08, -8.730431e-08, 
    -6.84361e-08, 1.349529e-07, -6.795915e-09, 2.031862e-08, -1.534312e-08, 
    4.798136e-08, 1.70175e-07, 1.401901e-07, -6.704278e-08, 9.163557e-09, 
    1.750719e-07, -3.715343e-09, 3.296662e-09, -5.849847e-08, 3.182939e-08, 
    -8.992612e-08, -4.634671e-08, -7.360258e-08, -2.314454e-08, 
    -3.257867e-09, -3.553794e-09, -6.286092e-08, -1.377619e-07, 4.429978e-09, 
    3.40921e-08, -5.394133e-08, 1.060482e-07, 2.773494e-07, -8.696077e-09, 
    2.601688e-07, 2.31438e-09, 7.927883e-09, -3.379167e-08, 1.345298e-07, 
    -1.722088e-08, -5.011297e-08, -1.903814e-07, -4.947573e-09, 9.115674e-09, 
    -2.197789e-08, 1.617292e-07, 4.19339e-08, -1.012012e-08, 1.057134e-08, 
    8.103086e-09, 4.958707e-08, 5.130119e-10, -4.882679e-09, -6.465768e-09, 
    -7.804545e-09, -7.488381e-09, -5.880918e-09, -2.269019e-09, -2.40032e-10, 
    -5.053664e-10, -3.714143e-08,
  1.174436e-08, -4.895526e-09, 2.434206e-09, 1.251789e-08, 8.98541e-09, 
    2.778978e-08, 2.879761e-08, 8.72916e-09, 2.177723e-08, 1.478901e-08, 
    2.223089e-09, -3.000594e-09, -2.641679e-08, 1.007714e-08, -1.266579e-08, 
    -1.508735e-08, -2.719051e-08, 4.108153e-08, -2.172922e-07, -5.677009e-09, 
    1.033059e-07, 2.658837e-07, 1.25386e-07, 1.428765e-08, -2.672039e-09, 
    -7.896682e-08, -3.621102e-08, -2.036239e-08, 4.522047e-08, -3.346344e-08, 
    -5.557814e-08, -1.502968e-08, 3.712955e-09, 7.10719e-09, -7.923478e-08, 
    5.144551e-08, -1.032072e-08, -3.357115e-09, -4.00442e-08, -3.940704e-08, 
    -5.889362e-09, 2.041759e-09, -1.419994e-08, -8.94839e-09, -3.47535e-09, 
    -3.977635e-08, 1.012174e-07, 8.999785e-08, 1.170755e-08, -5.933884e-10, 
    -1.527772e-08, -2.908149e-08, 1.284846e-07, -2.04718e-08, 5.975483e-08, 
    -2.001968e-09, -1.174794e-07, 2.284541e-07, 8.746232e-08, 2.874742e-09, 
    2.777313e-09, -1.085099e-07, -6.922409e-08, -8.437977e-08, -1.848827e-08, 
    8.068076e-08, -2.453879e-08, 2.84594e-08, -2.507119e-08, 4.645432e-08, 
    4.09176e-09, 1.947538e-07, -4.969519e-08, 1.033811e-09, 1.928777e-07, 
    -1.438337e-08, 2.600757e-09, -5.547219e-08, 3.358637e-08, 2.001951e-08, 
    -2.93075e-08, -6.089245e-08, -3.174029e-08, -4.23392e-08, -4.065271e-09, 
    -9.095953e-08, -1.818752e-07, 2.272719e-08, 3.896814e-08, -7.45481e-08, 
    6.339332e-08, 3.354541e-07, -8.164989e-09, 2.348796e-07, 4.348652e-08, 
    -1.316359e-07, -4.947902e-08, 5.72e-08, -2.085682e-08, -6.294505e-08, 
    -2.815393e-07, -4.078792e-08, 6.111726e-09, -1.974581e-08, 1.257026e-07, 
    3.968995e-08, 1.112255e-09, 1.616678e-08, 1.526172e-08, 6.224872e-08, 
    -2.078764e-10, -2.959666e-09, -8.679478e-09, -8.093537e-09, -8.60922e-09, 
    -4.684944e-09, -1.455504e-09, -3.147136e-10, -5.781757e-10, -3.589724e-08,
  5.021207e-09, -1.327714e-08, 1.626972e-09, -1.081946e-08, 1.218609e-09, 
    3.319826e-08, 3.114576e-08, 6.530513e-09, 3.112871e-08, -9.387122e-10, 
    -1.817114e-08, -4.727315e-08, -5.604159e-08, -4.416904e-08, 
    -1.419892e-08, -2.72551e-08, -2.631236e-08, 2.098091e-08, -2.154748e-07, 
    6.444691e-08, 3.545969e-07, 5.3897e-08, 1.816944e-07, 1.717865e-08, 
    -4.334345e-08, -1.017598e-07, -2.076092e-08, -1.256274e-08, 4.794094e-08, 
    -1.577234e-08, -6.688776e-08, -1.117303e-08, 1.41257e-08, 2.1451e-08, 
    -1.040549e-07, 1.318446e-07, -1.656299e-08, -8.282655e-10, -3.995831e-08, 
    -5.415975e-08, -1.463535e-07, 1.699277e-09, -1.432318e-08, -1.183189e-08, 
    7.77834e-09, -4.232277e-08, 9.439907e-08, 5.104363e-08, -1.709011e-08, 
    -3.148529e-09, -2.341466e-09, -1.37278e-08, 9.120083e-08, -1.87543e-08, 
    7.581212e-08, -5.012339e-09, -1.008153e-07, 1.395861e-07, 8.443988e-08, 
    -4.869719e-09, 1.660965e-10, -8.753352e-08, -7.950268e-08, -7.899546e-08, 
    -2.388726e-08, 6.362484e-09, -2.891909e-08, 5.354161e-08, -2.785043e-08, 
    4.546507e-08, 1.99347e-07, 2.649139e-07, -6.967946e-08, -4.963454e-09, 
    2.033775e-07, -2.540321e-08, 1.122316e-09, -3.752291e-08, 2.028578e-08, 
    -1.057139e-07, -1.150488e-08, -4.760007e-08, -1.627416e-08, 
    -7.905112e-08, 3.337971e-08, -1.141567e-07, -1.282596e-07, 4.421088e-08, 
    3.423046e-08, -9.968289e-09, 3.000821e-08, 3.470358e-07, -7.527717e-09, 
    2.289763e-07, 1.911261e-07, 1.487176e-08, -5.490148e-08, 3.620937e-08, 
    -2.555169e-08, -6.851226e-08, -2.046676e-07, -5.848264e-08, 6.218187e-09, 
    -1.65894e-08, 6.229163e-08, 1.340197e-08, -2.05215e-08, 1.328465e-08, 
    2.30765e-08, 6.117318e-08, -1.106059e-09, -1.197009e-09, -9.780138e-09, 
    -1.111414e-08, -3.736091e-09, -4.246931e-09, 2.414794e-09, -4.486935e-10, 
    -6.528893e-10, -3.023854e-08,
  -4.726417e-09, -3.176297e-08, 1.581839e-09, -3.416653e-08, -8.246161e-09, 
    2.921388e-08, 3.385708e-08, 1.111016e-08, 3.961804e-08, -6.911478e-09, 
    -2.186925e-08, -9.496762e-08, -2.435308e-08, -7.147037e-08, 4.444473e-09, 
    -3.297598e-08, -3.216021e-08, -1.067417e-08, -1.146394e-07, 1.322333e-07, 
    -1.443291e-07, -7.15404e-08, 2.563254e-07, 1.105459e-07, -7.780659e-08, 
    -6.914161e-08, -1.183207e-08, -2.001298e-08, 4.611547e-08, -1.56283e-08, 
    -7.23021e-08, -1.6988e-08, 6.294636e-08, -6.468758e-08, -1.106082e-07, 
    1.32366e-07, -1.93407e-08, -7.131575e-10, -2.688262e-08, -3.646248e-08, 
    -2.149865e-07, -6.423261e-08, -1.435978e-08, -7.196995e-09, -1.04933e-09, 
    -4.158414e-08, 1.287352e-07, 4.634001e-08, -3.055111e-08, -9.056947e-09, 
    1.008047e-08, -6.301661e-09, 5.011693e-08, -1.540611e-08, 8.995025e-08, 
    -3.351488e-09, -8.281427e-08, 1.778978e-07, 7.461817e-08, -2.362094e-08, 
    -2.748493e-09, -6.760365e-08, -5.488619e-08, -4.870235e-08, 
    -3.548939e-08, 1.983153e-09, -2.814636e-08, 9.023984e-08, -2.475963e-08, 
    3.996661e-08, 1.050148e-07, 1.925112e-07, -4.436583e-08, 5.218226e-10, 
    1.92079e-07, -3.103014e-08, 2.557726e-09, -2.46817e-08, 1.775634e-08, 
    -4.399658e-08, 2.652462e-08, -4.185155e-08, 1.028616e-08, -7.106519e-08, 
    7.201515e-08, -8.560687e-08, -1.391281e-07, 5.432139e-08, 3.76958e-08, 
    2.241813e-08, 1.134526e-08, 3.171186e-07, -6.533355e-09, 2.16013e-07, 
    4.983804e-08, 3.731957e-08, -4.397734e-08, -7.340168e-08, -3.061541e-08, 
    -6.721948e-08, -1.158926e-07, -5.174189e-08, 7.179295e-09, -1.258267e-08, 
    1.164358e-08, -1.058811e-08, -4.725007e-08, 4.08113e-09, 1.733724e-08, 
    4.310323e-08, -1.82381e-08, -1.228273e-09, -1.02757e-08, -1.722424e-08, 
    -1.168701e-09, -2.366278e-09, 8.072618e-09, -9.413839e-10, -7.121912e-10, 
    -5.139759e-08,
  -1.216063e-08, -5.439097e-08, 3.92879e-09, -2.036654e-08, -9.591758e-09, 
    2.773845e-08, 4.22931e-08, 1.777721e-08, 4.565936e-08, -2.342631e-09, 
    -1.915942e-08, -7.507833e-08, 8.636107e-09, -3.903369e-08, 1.509761e-08, 
    -4.196973e-08, -2.912736e-08, -1.03588e-08, -3.542112e-08, 6.557889e-08, 
    -8.725669e-08, -5.11468e-08, 1.547264e-07, 2.013846e-07, -2.296315e-08, 
    -3.662876e-08, 8.669986e-09, -6.874666e-08, 3.543232e-08, -1.012904e-08, 
    -6.132359e-08, -2.174761e-08, 5.104926e-08, -4.459343e-08, -8.859411e-08, 
    -4.747881e-08, -2.030699e-08, -2.847003e-10, -1.376202e-08, 
    -9.865771e-08, -2.412413e-07, 4.711867e-07, -1.941203e-10, 5.802388e-09, 
    -3.853984e-10, -4.139088e-08, 1.429248e-07, 4.892524e-08, -3.657474e-08, 
    -7.986813e-09, 2.239568e-08, -3.035757e-08, 6.363771e-08, -2.215866e-08, 
    9.116437e-08, -3.533728e-09, -6.155074e-08, 1.775081e-07, 4.165063e-08, 
    -5.698274e-08, -2.38856e-09, 6.486493e-08, -9.559722e-08, -1.129192e-08, 
    -3.196756e-08, -2.687784e-09, -2.326146e-08, 1.184517e-07, -2.772072e-08, 
    1.639228e-08, 2.779439e-08, 8.432221e-08, -2.922638e-08, 9.311179e-09, 
    1.473342e-07, -2.743263e-08, -2.421132e-09, -1.238959e-09, 8.065109e-09, 
    7.716062e-08, 8.117865e-08, -5.525897e-08, 3.286982e-08, -4.946787e-08, 
    -1.33432e-08, -7.606195e-08, -1.98675e-07, 4.354069e-08, 4.684767e-08, 
    4.331696e-09, 1.175795e-08, 2.886455e-07, -7.439837e-09, 1.808329e-07, 
    -4.846493e-08, 3.680921e-08, -1.610738e-08, -2.848719e-08, -3.26404e-08, 
    -7.570397e-08, -7.768449e-08, -3.607977e-08, 5.153666e-09, -5.705786e-09, 
    -2.191791e-08, -3.39719e-09, -1.605576e-08, 1.251465e-08, -3.524974e-09, 
    2.096249e-08, -4.365643e-08, -1.930857e-09, -8.763209e-09, -2.270008e-08, 
    -1.380977e-08, -7.315066e-10, 4.435464e-09, -2.080263e-09, -8.165273e-10, 
    -1.207713e-07,
  -9.053224e-09, -6.09574e-08, 2.789079e-09, 1.921023e-08, 3.281571e-09, 
    2.613058e-08, 5.130016e-08, 2.216518e-08, 5.345021e-08, 5.381673e-08, 
    -1.08256e-08, -2.396712e-08, 7.332289e-08, 3.758066e-08, 2.893705e-08, 
    -3.366324e-08, -2.720453e-08, 9.011501e-09, -2.932165e-08, 3.337266e-08, 
    7.310632e-09, -6.718585e-08, -3.425714e-08, 4.073058e-09, 1.025741e-07, 
    1.126421e-08, 2.133663e-08, -7.027154e-08, 3.216098e-08, -1.279284e-08, 
    -3.934963e-08, -1.635328e-08, 1.075239e-08, 2.169031e-09, -9.520215e-08, 
    8.356096e-09, -1.821343e-08, -1.212754e-09, -2.130685e-08, -1.144474e-07, 
    -2.421195e-07, 6.322955e-08, -3.833065e-08, 1.808859e-08, 5.347715e-09, 
    -2.899708e-08, 1.38597e-07, 6.681665e-08, -3.081452e-08, -3.877872e-09, 
    3.451331e-08, -8.072095e-08, 1.026929e-07, -2.38251e-08, 8.923804e-08, 
    -1.952685e-09, -4.976039e-08, 2.16808e-07, 5.87803e-08, -5.827374e-08, 
    3.785772e-11, 1.094469e-07, 1.572004e-07, 5.523248e-09, -9.788142e-09, 
    -1.34113e-08, -1.858314e-08, 2.881995e-08, -2.708441e-08, -2.970944e-08, 
    -2.772788e-08, 4.170749e-08, -3.269827e-08, 1.148317e-08, 1.011758e-07, 
    -1.669116e-08, -1.264513e-08, 9.494613e-09, 2.381733e-08, 2.227637e-08, 
    7.291965e-08, -8.396846e-08, 4.436799e-08, -2.373361e-08, -1.478668e-08, 
    -9.678945e-08, -2.712414e-07, 2.37643e-08, 5.588453e-08, -1.085664e-08, 
    -9.90633e-09, 2.623481e-07, -4.622336e-09, 1.204811e-07, -2.190279e-08, 
    2.760553e-08, 5.985605e-08, -1.824435e-08, -4.01966e-08, -9.333091e-08, 
    1.070254e-07, -8.519791e-09, 3.511715e-09, 1.771667e-09, -4.939204e-08, 
    -1.249759e-09, 1.165483e-08, 1.064075e-08, -2.52179e-08, 5.347033e-09, 
    -4.356878e-08, -1.031469e-08, -2.861384e-09, -2.810987e-08, -3.89947e-08, 
    -2.644811e-10, 2.329671e-09, -2.524544e-09, -9.586074e-10, -1.530628e-07,
  8.445227e-10, -3.411009e-08, -3.589491e-09, 3.678571e-08, 1.439281e-08, 
    1.40256e-08, 5.99278e-08, 1.911445e-08, 5.115709e-08, 9.110505e-08, 
    4.569466e-08, -3.464214e-08, -3.430836e-08, 5.325211e-08, -2.404585e-08, 
    -5.818383e-08, -1.408822e-08, 1.132111e-08, -6.056501e-08, 7.943129e-09, 
    4.898908e-08, -6.346107e-08, -1.671721e-07, -3.950998e-08, -6.383306e-08, 
    1.880342e-07, 2.206036e-09, -7.246234e-08, 3.154861e-08, -2.580595e-08, 
    -1.976167e-08, -7.774986e-09, 1.286372e-08, 9.203956e-08, -9.520835e-08, 
    1.552262e-07, -1.569075e-08, -3.916455e-09, -5.284204e-08, -4.930558e-08, 
    -1.968991e-07, -5.853957e-08, -4.728929e-08, 2.630704e-08, -6.247717e-09, 
    -1.744905e-08, 1.658603e-07, 1.066473e-07, -1.622806e-08, -2.424088e-10, 
    4.593204e-08, -1.113269e-07, 1.334269e-07, -2.842352e-08, 8.286473e-08, 
    -1.689443e-09, -4.621978e-08, 2.311104e-07, 1.249394e-08, -2.263266e-08, 
    -1.654001e-08, -2.663171e-09, 5.592761e-08, -3.445001e-08, -3.849652e-09, 
    -1.962661e-08, -7.955293e-09, -5.858908e-09, -1.662164e-08, 
    -5.709256e-08, -2.791188e-08, 7.403202e-08, -6.042455e-11, 6.341736e-09, 
    2.550299e-08, 6.441553e-09, -1.405675e-08, 1.60822e-08, 2.194731e-08, 
    -7.4355e-08, 5.149349e-08, -9.385369e-08, 8.801391e-08, -3.36683e-08, 
    8.547261e-09, 2.509371e-07, -2.266519e-07, 5.176673e-09, 6.238138e-08, 
    -2.0085e-08, 1.095908e-07, 2.305858e-07, -2.964782e-09, 6.851563e-08, 
    4.274744e-08, -4.110522e-08, 4.483505e-08, -4.614611e-08, -5.141573e-08, 
    -8.134774e-08, 3.956671e-08, -3.160152e-08, 2.472973e-09, 5.854716e-09, 
    -6.161525e-08, -1.883353e-08, 1.696532e-08, 1.089631e-09, -3.427539e-08, 
    -2.935337e-09, -3.330905e-08, -2.259293e-08, 1.684435e-08, -3.664076e-08, 
    -2.375089e-09, 5.916377e-10, 4.01991e-09, -2.103342e-09, -1.124747e-09, 
    -1.264636e-07,
  1.169764e-08, 3.071079e-09, -9.972666e-09, -2.244235e-09, -3.991829e-09, 
    -3.415721e-10, 4.403313e-08, -2.14946e-08, 4.730367e-08, 3.218287e-08, 
    -3.944598e-08, 6.498402e-08, 1.951227e-07, -1.092713e-07, -1.705718e-08, 
    -5.19907e-08, 6.316975e-09, 5.763638e-09, -8.011739e-09, -1.01839e-08, 
    1.847337e-08, -5.378621e-08, -1.491476e-07, -4.648479e-08, -1.121767e-07, 
    -9.121737e-08, -4.471588e-09, -7.065211e-08, 3.500321e-08, -1.752738e-08, 
    -5.977938e-09, -3.233993e-09, 2.127535e-07, 1.189291e-07, -7.488103e-08, 
    1.762514e-07, -1.431059e-08, -5.439119e-09, -7.168461e-08, -1.468955e-08, 
    -1.381771e-07, -7.523619e-08, 9.880461e-08, 2.971102e-09, 3.721397e-08, 
    -1.705763e-08, 2.06499e-07, 1.526067e-07, 2.917712e-08, 2.763372e-09, 
    5.569009e-08, -8.3609e-08, 1.590914e-07, -2.389362e-08, 7.280194e-08, 
    -2.742411e-09, -4.473242e-08, 2.256295e-07, 6.060701e-08, -3.771757e-08, 
    -5.647342e-07, -1.605582e-08, 9.916943e-08, -2.974609e-08, -1.574109e-08, 
    -1.45854e-08, -3.751722e-09, 5.332521e-08, -2.3415e-08, -5.473663e-08, 
    -3.627594e-08, 1.08414e-07, 7.494913e-08, 5.792702e-08, 5.785342e-08, 
    1.862662e-08, -5.593193e-09, 2.523132e-08, 2.14311e-08, -3.14306e-08, 
    4.650934e-08, -7.660979e-08, 8.397666e-08, -4.812165e-08, 1.201537e-07, 
    2.375618e-07, -1.564104e-07, -5.983622e-09, 6.904695e-08, -3.949123e-08, 
    -5.947624e-08, 2.15332e-07, -4.011611e-09, 7.081975e-08, 3.993313e-08, 
    -1.490985e-07, 2.562896e-08, 2.639524e-09, -6.363331e-08, -9.582546e-08, 
    -6.972874e-08, 1.751743e-07, 4.945093e-09, 7.553638e-09, -4.859027e-08, 
    -4.097393e-08, 1.436268e-08, -6.245784e-09, -3.013935e-08, -5.559343e-09, 
    -2.842495e-08, -2.452867e-08, 1.467737e-08, -4.233772e-08, 3.098364e-09, 
    5.035304e-10, 6.556775e-09, -2.358739e-09, -1.118565e-09, 8.589603e-08,
  1.395335e-08, 4.809851e-08, -2.058243e-08, -1.801993e-08, 8.3445e-09, 
    -4.695869e-08, -3.590799e-09, -5.483992e-08, 1.320392e-07, -2.562899e-08, 
    -2.339073e-08, -1.690216e-08, 1.172772e-07, -1.155271e-07, 1.181755e-07, 
    2.516366e-09, 2.087438e-08, 1.289141e-08, 2.343083e-08, -8.323127e-09, 
    8.309712e-09, -3.14559e-08, -1.27275e-07, 2.071909e-08, -1.929101e-07, 
    -6.718108e-08, -3.788614e-09, -6.347284e-08, 4.010724e-08, 5.214474e-09, 
    1.101512e-09, -6.618052e-09, 1.630225e-07, 5.106824e-08, -4.828155e-08, 
    1.426528e-07, -1.600492e-08, -2.582993e-09, -4.057654e-08, 7.564815e-09, 
    -1.244923e-07, -3.497215e-07, -3.246606e-08, -1.048217e-08, 1.699607e-08, 
    -1.966885e-08, 3.049687e-07, 1.991967e-07, 3.067692e-08, 3.490115e-09, 
    6.27617e-08, 6.04922e-08, 1.777268e-07, -1.035385e-08, 5.819322e-08, 
    -2.997922e-09, -4.109972e-08, 1.710289e-07, 1.294144e-07, -3.558299e-08, 
    1.634509e-07, -1.114779e-08, -8.874281e-09, -1.333444e-08, -2.000136e-08, 
    -2.744457e-08, -2.579441e-09, 2.175545e-08, -5.158938e-08, -5.505797e-08, 
    -2.342938e-08, 1.187567e-07, 5.833738e-08, 3.419893e-08, 6.982199e-08, 
    -1.593946e-08, -3.819423e-09, 2.799504e-08, 2.146891e-08, -1.167029e-08, 
    7.813981e-08, -4.193269e-08, 7.229175e-08, 4.089202e-09, 6.692233e-08, 
    -5.850666e-09, -7.855704e-08, -1.603109e-08, 3.950812e-08, -1.212129e-08, 
    -7.362098e-08, 1.97558e-07, -5.647621e-09, 6.631057e-09, 6.685434e-08, 
    3.30806e-09, -1.403521e-08, 2.252034e-08, -5.894947e-08, -1.307347e-07, 
    -1.053905e-07, -4.670363e-08, 9.515254e-08, 8.303147e-09, -2.156742e-08, 
    -4.171318e-08, 2.569107e-08, -9.245582e-09, -2.135869e-08, -4.508479e-09, 
    -2.661238e-08, -2.001559e-08, -3.968808e-10, -3.281559e-08, 3.868649e-09, 
    -1.881744e-10, 8.658617e-09, -2.683407e-09, -1.074795e-09, 6.193557e-08,
  -3.503385e-08, 2.936883e-08, -7.307312e-08, 5.167078e-08, 5.41155e-08, 
    -1.168559e-07, -1.477679e-08, -4.408037e-08, 1.98031e-07, -4.855451e-09, 
    -3.300556e-09, -3.22616e-08, 1.173862e-08, 8.696145e-08, 4.831088e-08, 
    1.96241e-08, 4.370973e-08, 3.552958e-08, -7.108723e-08, 5.279094e-08, 
    6.624532e-10, -1.469834e-08, -5.763673e-08, 8.597453e-09, -9.825146e-08, 
    2.81625e-09, 3.18596e-09, -5.693414e-08, 4.447804e-08, 6.785172e-09, 
    6.950131e-09, -3.216201e-10, 8.484903e-08, 1.337479e-07, 1.938452e-08, 
    -4.168589e-08, -4.200148e-08, 6.008307e-09, -2.382092e-08, 3.084938e-08, 
    -8.581199e-08, -3.359228e-07, -4.230782e-08, 4.102784e-09, -9.310952e-11, 
    -1.74806e-08, 3.743066e-07, 2.340787e-07, 2.970337e-08, 2.705548e-09, 
    6.732385e-08, 1.17618e-07, 1.633537e-07, -1.264539e-09, 3.494734e-08, 
    -1.938872e-09, -3.825744e-08, 8.714137e-08, 1.236144e-07, -3.334405e-08, 
    -1.94105e-07, -2.280001e-08, -1.310252e-08, -1.629228e-08, -1.714193e-08, 
    -7.379526e-09, 6.223217e-10, 1.771184e-08, -4.133301e-08, -2.636875e-08, 
    -2.816842e-08, 1.026182e-07, 2.353318e-10, -1.980027e-08, 6.326347e-08, 
    -2.564093e-08, -6.058798e-10, 3.456873e-08, 1.595734e-08, 1.867079e-09, 
    1.12868e-07, 1.690287e-08, 6.323705e-08, 4.726244e-07, 4.057893e-08, 
    -2.355785e-07, -1.108749e-07, -3.209846e-08, 9.866291e-09, 5.472145e-09, 
    1.674607e-08, 1.752102e-07, -6.163646e-09, -2.14824e-08, 1.235499e-07, 
    1.673925e-09, 8.881898e-09, 7.133963e-09, -5.043387e-08, -8.946124e-08, 
    -7.800952e-08, -3.60284e-08, 1.392698e-07, 7.997919e-09, 3.430716e-08, 
    -1.009147e-07, 6.607002e-08, -1.631236e-08, -1.521414e-08, -2.359116e-09, 
    -2.569152e-08, -1.722913e-08, -6.297569e-09, -1.043122e-08, 3.942546e-09, 
    -5.194692e-10, 9.026522e-09, -2.469605e-09, -1.064031e-09, 5.505808e-08,
  -1.983512e-07, -3.465378e-07, -1.903831e-07, 2.33635e-07, 1.804526e-07, 
    -1.146879e-07, 1.028459e-07, -2.955125e-08, 1.268137e-08, -1.420716e-08, 
    1.223219e-08, -2.695839e-08, -4.514521e-08, 8.981948e-08, 1.550263e-07, 
    2.885698e-08, 3.021861e-08, 2.930551e-08, -1.10541e-07, 1.93849e-07, 
    4.405473e-08, -1.97413e-07, 3.313534e-08, 6.320704e-09, -5.971458e-09, 
    3.136921e-08, -8.090126e-09, -5.578528e-08, 6.564943e-08, -1.891334e-08, 
    9.22131e-09, 1.219024e-08, 1.793097e-08, 1.012272e-07, 2.359332e-07, 
    -7.190073e-08, -3.789707e-08, 1.861397e-08, -5.278764e-09, 4.829652e-08, 
    -8.931906e-09, -1.107322e-07, -2.147351e-08, -2.692726e-08, 
    -1.649602e-08, -1.713573e-08, 4.103559e-07, 2.381371e-07, 6.178792e-08, 
    2.338886e-09, 7.016733e-08, 1.814275e-07, 1.006226e-07, 2.554622e-08, 
    1.26757e-08, -3.151513e-09, -4.860823e-08, 6.482346e-08, -5.820027e-09, 
    -3.336409e-08, 3.207634e-08, 8.494112e-10, -1.225101e-07, -3.984668e-08, 
    -3.041708e-08, -1.043719e-08, 3.822436e-09, 7.237475e-09, 3.194526e-08, 
    6.109246e-09, -1.864083e-08, 8.307944e-08, -1.138329e-08, -2.959513e-08, 
    6.623758e-08, -2.465464e-08, -2.27799e-08, 3.397201e-08, 1.220969e-08, 
    4.165878e-08, 5.692846e-08, 5.568662e-08, 4.345054e-08, 1.791612e-07, 
    4.474992e-08, -6.34289e-08, -3.110091e-08, -6.122644e-08, -8.986991e-09, 
    8.081201e-09, 1.982478e-07, 1.100718e-07, -2.276835e-09, -1.744906e-08, 
    2.657833e-08, 1.860041e-09, 5.337085e-09, -5.201912e-09, -2.713472e-08, 
    -2.364199e-08, -6.181779e-09, -7.996636e-08, 1.634826e-07, 6.644193e-09, 
    6.078488e-08, -2.84918e-08, 1.098197e-07, -1.990492e-08, -1.247992e-08, 
    -9.395649e-10, -2.50979e-08, -1.603229e-08, -6.292566e-11, -2.5031e-09, 
    3.684875e-09, -6.629307e-10, 8.63453e-09, -2.377664e-09, -8.150352e-10, 
    1.769655e-08,
  -3.0835e-07, -8.87913e-07, -1.009169e-07, 2.075123e-07, 3.57908e-07, 
    1.467196e-07, 8.954913e-08, 8.642138e-08, -4.862756e-08, -2.010955e-08, 
    1.903078e-08, -2.228734e-08, -2.673862e-07, 7.169621e-08, -4.411453e-08, 
    3.353504e-08, 3.505533e-08, 1.358501e-08, -1.30711e-07, 1.794149e-09, 
    -2.346457e-08, -5.42488e-08, 7.621736e-09, 8.579889e-09, 1.746531e-08, 
    1.784639e-08, 7.18382e-08, -5.863905e-08, 9.26637e-08, -4.068505e-08, 
    -1.203415e-08, 4.075275e-09, -8.601745e-08, 2.926268e-07, 1.425498e-07, 
    -1.172651e-08, -2.048127e-08, 2.68203e-08, 5.821846e-09, 5.966774e-08, 
    6.966737e-09, -1.097879e-08, -1.525734e-08, -1.921701e-08, 8.917539e-09, 
    1.797918e-08, 4.279886e-07, 2.150607e-07, 5.764224e-08, 2.115982e-09, 
    7.018102e-08, 8.467003e-08, 8.366339e-08, 4.663656e-08, 1.645887e-09, 
    -5.269783e-09, -5.796636e-08, 3.80695e-08, 6.499477e-10, -3.076408e-08, 
    1.549603e-08, 1.067195e-08, -5.994735e-08, -4.401508e-08, -2.793075e-08, 
    -9.681287e-09, 1.953424e-09, 1.57242e-08, 5.978114e-08, 7.597066e-09, 
    -2.496512e-08, 6.301337e-08, 1.128342e-10, -2.861185e-08, 7.266269e-08, 
    -2.94595e-08, -4.163198e-08, 4.204162e-08, 4.486893e-09, 9.75835e-08, 
    -1.943238e-08, 6.09496e-08, 3.729605e-08, -1.733956e-07, -4.991591e-09, 
    6.394094e-08, -2.820053e-08, -9.744082e-08, -1.650657e-08, 7.830238e-09, 
    1.734264e-08, 8.798287e-08, -6.841617e-09, -2.08662e-09, 4.495803e-09, 
    4.086383e-09, -1.848485e-08, 6.295011e-09, -6.247564e-08, -2.724036e-08, 
    -3.928818e-08, -6.261651e-08, 2.800473e-08, 6.695544e-09, -7.861388e-09, 
    -1.934319e-08, 1.586981e-07, -2.200665e-08, -1.039024e-08, 3.087337e-09, 
    -2.469409e-08, -1.489337e-08, 3.147022e-09, -1.664091e-09, 3.081198e-09, 
    -4.293725e-10, 6.103591e-09, -2.422109e-09, -8.463914e-10, 1.083157e-08,
  -1.825368e-07, -6.295523e-07, 1.082062e-07, 3.438157e-08, -9.591628e-08, 
    9.995046e-08, 1.316059e-07, 5.876194e-08, -2.239409e-08, -1.977156e-08, 
    -5.60027e-09, -2.106901e-09, -8.667104e-08, 1.030611e-08, -1.199811e-08, 
    2.331777e-08, 7.22423e-10, -9.429471e-09, -1.590652e-08, -1.14224e-08, 
    -1.64319e-08, 6.697917e-09, 8.335462e-09, 8.880704e-09, 3.456574e-08, 
    1.320808e-08, 6.688305e-08, -5.769522e-08, 2.919177e-08, -6.645524e-08, 
    -7.160753e-08, -5.548219e-08, -9.293768e-08, 1.856401e-07, -5.708728e-09, 
    4.621637e-08, -1.484715e-08, 3.140778e-08, -2.896837e-08, 6.784759e-08, 
    -3.436272e-08, 1.752477e-08, -1.167018e-08, -2.0018e-08, -2.77135e-08, 
    8.495175e-08, 4.79133e-07, 1.943907e-07, 3.131844e-08, 1.786645e-09, 
    8.387215e-08, 1.885098e-09, 6.900513e-08, 3.228187e-08, -3.511383e-09, 
    -2.353602e-09, -4.141117e-08, 4.027594e-08, 1.833826e-09, -1.68759e-08, 
    1.712777e-08, 1.16824e-08, 4.017863e-09, -5.508174e-08, -3.631936e-08, 
    -9.180951e-09, -1.738869e-08, -6.237372e-09, 5.970531e-08, 2.419159e-08, 
    -3.843007e-08, 4.450538e-08, -1.84728e-08, 3.549911e-08, 7.550631e-08, 
    -3.093356e-08, 5.069353e-09, 2.586108e-08, 5.582415e-10, 2.228232e-07, 
    -9.484307e-08, 4.655379e-08, 2.98424e-08, -8.215449e-08, 2.444665e-09, 
    1.634903e-07, -1.339987e-08, -8.927424e-08, -2.835519e-08, 2.08118e-08, 
    -1.569384e-08, 8.016453e-08, -2.867353e-09, 9.050393e-09, 5.681085e-08, 
    1.003201e-08, -4.286022e-08, 6.491194e-08, -5.388966e-08, 1.288976e-08, 
    -3.687097e-08, 9.611554e-09, -3.744179e-08, 6.960462e-09, -1.430975e-07, 
    -4.396753e-08, 1.853302e-07, -2.145299e-08, 2.884804e-10, 7.935057e-09, 
    -2.432972e-08, -1.400764e-08, 3.407138e-09, -1.699902e-09, 2.732975e-09, 
    6.11692e-10, 9.655139e-09, -1.916298e-09, -1.127475e-09, -1.548472e-09,
  -1.195431e-07, 2.373156e-08, 1.072569e-07, 4.576123e-08, -5.073537e-08, 
    1.603894e-08, -2.661943e-08, -5.369316e-09, -9.446921e-09, -7.139988e-09, 
    -5.402853e-09, -3.135028e-09, 1.398769e-08, 1.713931e-08, -1.551791e-08, 
    2.343901e-08, -1.141788e-08, -2.984825e-08, 2.816478e-09, -1.432488e-08, 
    -1.133913e-08, 4.654714e-08, 7.17273e-09, 9.138489e-09, 4.093863e-08, 
    1.042019e-08, 6.06035e-08, -3.952482e-08, -1.021601e-08, -6.167454e-08, 
    -1.040775e-07, 3.618925e-08, -1.105938e-07, 2.01741e-07, -4.616481e-09, 
    1.01829e-07, -1.395681e-08, 3.219907e-08, -4.000549e-08, 7.30218e-08, 
    -9.316072e-08, 3.060575e-08, -1.106355e-08, -2.271646e-09, 9.19124e-09, 
    2.032277e-08, 5.201671e-07, 1.850526e-07, 6.488676e-09, 9.378169e-10, 
    8.325428e-08, -6.080882e-09, 4.951398e-08, 2.869251e-08, -7.709562e-09, 
    -1.575984e-09, -8.497636e-09, 4.494022e-08, 1.227356e-10, 9.543655e-09, 
    2.004776e-08, 1.199203e-08, 2.296838e-08, -5.639806e-08, 5.818742e-09, 
    4.809533e-08, -3.629395e-08, -2.52453e-09, 1.001649e-08, -1.851686e-08, 
    -3.964715e-09, 2.098625e-08, -1.020192e-08, 1.113824e-08, 7.419501e-08, 
    -3.265234e-08, 1.833567e-08, 1.899156e-08, -2.103713e-09, 1.066783e-07, 
    -3.571733e-08, 4.5442e-08, 4.462453e-08, -3.809214e-08, 2.678667e-08, 
    7.110339e-08, -1.477508e-08, -2.064507e-08, -2.420759e-08, 3.658289e-08, 
    -2.641184e-08, 6.99061e-08, -6.69246e-10, 1.440053e-08, 1.201684e-07, 
    1.979763e-08, -4.660706e-08, 1.729283e-07, -5.551726e-08, -1.968672e-08, 
    -7.282915e-08, 2.463717e-08, -4.446692e-08, 7.732858e-09, -2.814878e-07, 
    -6.881464e-09, 2.016922e-07, -1.986473e-08, 5.101356e-09, 1.549984e-08, 
    -2.394245e-08, -1.323758e-08, 3.279638e-09, -1.655394e-09, 1.294779e-09, 
    -5.24119e-10, 7.43816e-09, -1.751975e-09, -1.240124e-09, -1.529997e-09,
  -1.324642e-07, 1.760009e-08, 1.019365e-07, 4.620426e-08, -2.433001e-08, 
    -1.013746e-09, -2.731565e-08, -1.019657e-08, -6.200821e-09, 
    -2.267825e-09, -5.496645e-09, -3.908553e-09, 1.233809e-08, 1.216233e-08, 
    -1.675483e-08, 2.121954e-08, -1.806433e-08, 9.555663e-09, -1.484869e-08, 
    -1.547085e-08, -9.161113e-09, 5.278264e-08, 4.20539e-09, 8.992515e-09, 
    4.413539e-08, 1.047135e-08, 6.455355e-08, 2.884724e-08, -9.152814e-09, 
    -8.130382e-08, -1.095575e-07, -5.285949e-08, -1.8432e-07, 2.298167e-07, 
    -3.869786e-09, 1.756162e-07, -1.485591e-08, 2.777549e-08, -6.70093e-09, 
    7.423299e-08, -9.348246e-08, 3.503362e-08, -1.218115e-08, -2.499174e-10, 
    2.519062e-08, -3.382638e-09, 5.334191e-07, 1.850331e-07, 2.237199e-09, 
    1.021426e-09, 8.0487e-08, -9.838118e-09, 3.340084e-08, 2.856487e-08, 
    -1.003582e-08, -3.878995e-10, 8.164307e-09, 3.422135e-08, 8.550829e-09, 
    2.596212e-08, 2.151944e-08, 1.244575e-08, 2.122999e-08, -4.813432e-08, 
    2.202578e-08, 4.427989e-08, 7.00735e-08, -6.739208e-08, 2.40924e-08, 
    -3.864591e-08, 9.976134e-09, 3.005312e-09, -7.483209e-09, 1.743365e-08, 
    7.045324e-08, -2.66898e-08, 3.935183e-08, 5.972822e-09, -3.767155e-09, 
    5.72918e-08, -3.385099e-08, 4.537283e-08, 5.121211e-08, -1.381397e-08, 
    -5.264974e-08, 5.620529e-08, -1.462024e-08, 5.247398e-08, -2.00609e-08, 
    4.270169e-08, -3.09135e-08, 6.984713e-08, -1.880096e-10, 1.454673e-08, 
    -3.51713e-08, 2.846615e-08, -4.18383e-08, 4.019148e-08, -6.48073e-08, 
    -5.565127e-09, -5.308493e-09, 3.264868e-08, -3.982266e-08, 8.187207e-09, 
    -2.87468e-07, 3.654725e-08, 1.982091e-07, -2.27426e-08, 5.85942e-09, 
    1.372905e-08, -2.359661e-08, -1.285787e-08, 3.259402e-09, -1.530907e-09, 
    -3.274181e-11, 2.007857e-09, 7.891401e-09, -1.579828e-09, -3.122366e-09, 
    -1.711896e-09,
  -7.704892e-08, 2.280143e-08, 1.059072e-07, 4.485906e-08, -1.321467e-08, 
    -6.293533e-09, -3.060887e-08, -1.138216e-08, 2.785328e-12, -8.525944e-10, 
    -5.742834e-09, -4.584592e-09, 9.309076e-09, 8.432096e-09, -1.594952e-08, 
    2.463662e-08, -6.83923e-09, 6.371181e-09, -1.653355e-08, -1.595635e-08, 
    -8.181871e-09, 6.067791e-08, 5.33845e-09, 9.341363e-09, 4.689497e-08, 
    8.214386e-09, 1.642337e-08, 1.145776e-08, -8.835798e-09, -1.061237e-07, 
    -8.014825e-08, -6.210922e-08, -3.346502e-07, 2.379144e-07, -2.784702e-09, 
    2.398991e-07, -1.637741e-08, 1.514597e-08, -3.680555e-09, 7.392484e-08, 
    -9.880252e-08, 3.782458e-08, -1.278241e-08, -8.048218e-09, 1.783354e-08, 
    -1.349605e-08, 5.017925e-07, 1.924582e-07, -4.66099e-09, 4.363159e-10, 
    7.712397e-08, -1.186851e-08, 2.32909e-08, 3.226138e-08, -7.406578e-09, 
    -2.145043e-09, -2.43989e-09, 3.186809e-08, 3.6747e-09, 7.854311e-09, 
    2.165945e-08, 1.192853e-08, 1.557004e-08, -4.032346e-08, 3.637134e-08, 
    1.903135e-08, -2.737266e-08, -3.438123e-08, -1.149607e-08, 4.791565e-08, 
    1.028354e-09, -4.743299e-09, -6.102994e-09, 1.940219e-08, 6.448304e-08, 
    -2.862481e-08, 5.412792e-08, 1.968658e-09, 7.485967e-10, 5.702526e-08, 
    -3.837988e-08, 3.471851e-08, 5.022287e-08, -8.340635e-10, -5.420878e-08, 
    5.826081e-08, -1.452412e-08, 5.151747e-08, -1.941332e-08, 4.688974e-08, 
    -3.258361e-08, 6.462168e-08, 1.346024e-09, 1.217832e-08, -3.65049e-08, 
    3.559016e-08, -4.025184e-08, 3.801148e-08, -4.620091e-08, -2.49662e-09, 
    5.426671e-09, 3.650581e-08, -9.455309e-08, 8.483298e-09, -1.027285e-07, 
    -2.065184e-08, 1.846381e-07, -2.736743e-08, 4.568562e-09, 1.115274e-08, 
    -2.114501e-08, -1.234645e-08, 3.124057e-09, -1.477645e-09, -5.590493e-09, 
    4.39494e-09, 8.751414e-09, -1.366981e-09, -4.561215e-09, -1.414776e-09,
  -6.315184e-08, 2.2336e-08, 1.071549e-07, 4.620375e-08, -9.209941e-09, 
    -8.088307e-09, -3.128815e-08, -1.16259e-08, -1.297735e-10, -6.085088e-10, 
    -6.041603e-09, -5.168829e-09, 7.867641e-09, 6.12755e-09, -1.674374e-08, 
    2.968787e-08, 1.174317e-09, -5.072309e-09, -2.075105e-08, -1.688767e-08, 
    -7.558185e-09, 6.590773e-08, 7.583537e-09, 9.795087e-09, 4.693919e-08, 
    5.801496e-09, 2.238568e-08, -2.897974e-08, -8.911172e-09, -1.684327e-09, 
    -1.427753e-08, -1.245441e-07, -3.629934e-07, 2.072482e-07, -1.678757e-09, 
    2.69462e-07, -1.814936e-08, 2.956682e-09, 1.941504e-08, 7.245437e-08, 
    -9.982819e-08, 3.878637e-08, -1.257123e-08, -6.083146e-09, -2.985587e-09, 
    -1.756865e-08, 4.578425e-07, 2.052606e-07, -8.366135e-09, -2.989253e-11, 
    7.649024e-08, -1.319148e-08, 1.69886e-08, 3.153865e-08, -1.359792e-08, 
    9.472387e-10, -1.775066e-08, 2.502888e-08, 1.344847e-09, 3.016879e-09, 
    2.117002e-08, 1.078428e-08, 1.33486e-08, -5.12607e-08, 2.707499e-08, 
    1.754034e-08, -4.210591e-08, -3.446274e-08, 2.25387e-08, 6.058707e-08, 
    -2.516856e-09, -1.188533e-08, -5.410982e-09, 2.007022e-08, 5.910849e-08, 
    -1.043196e-08, 5.264238e-08, 1.114282e-08, -2.743432e-10, 5.222176e-08, 
    -4.028834e-08, 2.696819e-08, 4.352717e-08, 6.047173e-09, -5.965109e-08, 
    6.066949e-08, -1.365089e-08, 4.942359e-08, -2.126227e-08, 4.839114e-08, 
    -3.269128e-08, 5.956789e-08, 2.663171e-09, 7.295535e-09, -8.409927e-09, 
    4.189052e-08, -3.973583e-08, 4.049554e-08, -3.699364e-08, -4.945946e-10, 
    1.391908e-08, 3.912028e-08, -8.953675e-08, 7.99222e-09, -6.97093e-08, 
    -2.700693e-08, 2.019025e-07, -3.346048e-08, 2.450804e-09, 8.651284e-09, 
    -1.818199e-08, -1.095628e-08, 3.044818e-09, -1.236856e-09, -2.873668e-08, 
    2.888828e-09, 2.751989e-09, -8.662617e-10, -9.598793e-10, 3.632863e-10,
  -4.991779e-08, 2.063911e-08, 1.060442e-07, 4.404814e-08, -8.066365e-09, 
    -8.626728e-09, -3.117458e-08, -1.152881e-08, -1.23481e-09, -6.115783e-10, 
    -6.40938e-09, -2.202739e-09, 7.301594e-09, 7.362758e-09, -1.640007e-08, 
    3.117277e-08, -1.3957e-09, -6.894084e-09, -2.368563e-08, -1.744246e-08, 
    -7.130382e-09, 6.884619e-08, 8.646737e-09, 1.000654e-08, 4.566317e-08, 
    5.419736e-09, 2.00892e-08, -3.527401e-08, -9.145481e-09, 4.177542e-08, 
    1.786356e-08, -4.560144e-08, -4.054534e-07, 2.187679e-07, -7.416361e-10, 
    3.044624e-07, -1.994524e-08, 6.45862e-09, 9.155031e-09, 7.02552e-08, 
    -9.906854e-08, 3.974191e-08, -1.22883e-08, -1.047114e-08, -8.010545e-09, 
    -2.04073e-08, 3.969558e-07, 2.205403e-07, -1.002278e-08, -7.378418e-10, 
    7.74658e-08, -1.451969e-08, 1.512955e-08, 3.281626e-08, -1.387639e-08, 
    -1.481169e-09, -3.036445e-08, 1.822897e-08, -1.866806e-09, -2.067608e-09, 
    2.015196e-08, 1.037421e-08, 1.223844e-08, -7.045978e-08, 2.866847e-08, 
    4.004295e-08, -2.446603e-08, -7.277396e-08, 1.702693e-08, 3.677422e-08, 
    -3.809515e-08, -6.392781e-09, -5.142681e-09, 2.031999e-08, 5.314228e-08, 
    -4.413039e-09, 5.250341e-08, 6.744699e-09, -2.251147e-09, 4.927421e-08, 
    -3.972434e-08, 2.14539e-08, 4.39249e-08, 9.315215e-09, -6.209081e-08, 
    6.179806e-08, -1.292761e-08, 4.740713e-08, -2.132357e-08, 4.728651e-08, 
    -3.241252e-08, 5.567253e-08, 3.477311e-09, 4.263098e-09, -5.797745e-09, 
    4.689461e-08, -4.001871e-08, 3.969257e-08, -3.469319e-08, -5.226291e-10, 
    1.589075e-08, 4.144464e-08, -9.032268e-08, 7.088424e-09, -8.248372e-08, 
    -2.797509e-08, 3.885573e-07, -3.738609e-08, 6.32042e-10, 5.647905e-09, 
    -1.521067e-08, -8.386621e-09, 3.200682e-09, -8.289476e-10, -3.950487e-08, 
    1.098272e-09, -3.777814e-10, -2.878501e-09, 4.475268e-09, 1.321439e-09,
  -4.377569e-08, 1.876606e-08, 1.015079e-07, 4.090975e-08, -8.288566e-09, 
    -9.070391e-09, -3.047262e-08, -1.121236e-08, -3.104105e-09, 
    -8.557208e-10, -7.020617e-09, -2.16869e-09, 6.790856e-09, 1.056731e-08, 
    -1.621072e-08, 3.191559e-08, -5.798596e-10, -8.111556e-09, -2.557412e-08, 
    -1.817614e-08, -6.911932e-09, 7.101346e-08, 9.298333e-09, 1.016883e-08, 
    4.345748e-08, 4.363756e-09, 1.881983e-08, -4.303399e-08, -9.527184e-09, 
    1.558908e-08, 3.969728e-08, -3.955381e-08, -4.502925e-07, 2.386647e-07, 
    1.367653e-10, 3.238476e-07, -2.152539e-08, 6.866372e-09, -2.85786e-09, 
    6.82808e-08, -9.738564e-08, 3.871537e-08, -1.204816e-08, -1.10698e-08, 
    -1.582453e-08, -2.474417e-08, 3.525229e-07, 2.390771e-07, -1.178155e-08, 
    -1.860315e-09, 7.811833e-08, -1.584408e-08, 1.349691e-08, 2.796726e-08, 
    1.947868e-09, -1.942965e-09, -3.98926e-08, 1.098954e-08, -6.005506e-09, 
    -5.725738e-09, 1.849946e-08, 1.015371e-08, 1.201579e-08, -1.085677e-07, 
    3.163164e-08, 4.953631e-08, -1.730336e-08, -8.928782e-08, 1.827289e-08, 
    3.212028e-08, -4.576179e-08, -4.857225e-08, -4.588742e-09, 1.986268e-08, 
    4.675075e-08, -3.062382e-09, 5.193729e-08, 3.699341e-09, -2.917133e-09, 
    4.692458e-08, -3.807446e-08, 1.668974e-08, 4.321316e-08, 1.034346e-08, 
    -6.148287e-08, 6.048776e-08, -1.162061e-08, 4.511298e-08, -2.077393e-08, 
    4.586445e-08, -3.219134e-08, 5.384686e-08, 3.598473e-09, -6.778134e-10, 
    1.103786e-09, 5.079158e-08, -3.889297e-08, 3.831292e-08, -3.346133e-08, 
    -1.4021e-09, 2.140234e-08, 4.310219e-08, -9.045206e-08, 5.934822e-09, 
    -8.941117e-08, -2.813476e-08, 4.579215e-07, -3.904108e-08, -2.961542e-10, 
    3.108767e-09, -1.443118e-08, -4.887283e-09, 4.167532e-09, -5.733227e-10, 
    -4.953006e-08, -9.195106e-10, -4.267676e-09, -1.981846e-10, 4.359947e-09, 
    2.770548e-10,
  -4.44856e-08, 1.633049e-08, 9.645811e-08, 3.8324e-08, -9.036228e-09, 
    -9.613643e-09, -2.915743e-08, -1.070913e-08, -3.576872e-09, -1.7057e-09, 
    -7.819892e-09, -1.969227e-09, 5.637901e-09, 1.112716e-08, -1.584141e-08, 
    2.388283e-08, 1.161811e-09, -9.291966e-09, -2.707976e-08, -1.917016e-08, 
    -7.217693e-09, 7.228488e-08, 9.92992e-09, 1.037944e-08, 4.185682e-08, 
    2.585296e-09, 1.890027e-08, -4.231862e-08, -1.009431e-08, -4.872447e-09, 
    5.021462e-08, -3.801284e-08, -4.922148e-07, 2.845799e-07, 1.247656e-09, 
    3.319013e-07, -2.273805e-08, 5.91244e-09, -1.235918e-08, 5.892052e-08, 
    -9.614899e-08, 3.662336e-08, -1.182806e-08, -1.025685e-08, -1.876396e-08, 
    -2.86272e-08, 2.836142e-07, 2.608166e-07, -1.359862e-08, -8.561386e-09, 
    8.37926e-08, -1.737766e-08, 1.237017e-08, 2.847752e-08, 2.13019e-08, 
    -4.147296e-09, -4.470581e-08, 3.081301e-09, -1.06838e-08, -8.091789e-09, 
    1.578616e-08, 9.597954e-09, 1.255711e-08, -1.820987e-07, 2.306482e-08, 
    5.768965e-08, -1.472807e-08, -1.032482e-07, 2.244354e-08, 2.206099e-08, 
    -4.804241e-08, -7.727482e-08, -3.767184e-09, 1.876077e-08, 4.031127e-08, 
    -2.275971e-08, 5.033613e-08, 2.241876e-09, -2.283505e-09, 4.551924e-08, 
    -3.669174e-08, 1.335026e-08, 4.109773e-08, 9.963003e-09, -5.964381e-08, 
    5.97426e-08, -1.017685e-08, 4.18874e-08, -2.275611e-08, 5.099866e-08, 
    -3.142583e-08, 5.219841e-08, 3.298652e-09, -4.145774e-09, 6.963944e-09, 
    5.393553e-08, -3.957667e-08, 3.868394e-08, -3.127974e-08, -1.443244e-09, 
    2.563701e-08, 4.438503e-08, -9.262362e-08, 4.849014e-09, -1.027285e-07, 
    -2.768974e-08, -3.883957e-08, -3.943848e-08, -6.635332e-10, 1.611568e-09, 
    -1.464656e-08, -1.839624e-09, 4.663264e-09, -9.053451e-10, -5.290536e-08, 
    -4.270873e-10, -1.041626e-08, -3.053078e-09, -1.499814e-10, -8.100187e-11,
  -4.502635e-08, 1.158708e-08, 9.177359e-08, 3.57777e-08, -1.037017e-08, 
    -1.062676e-08, -2.60452e-08, -9.512632e-09, -1.868329e-09, -3.99973e-09, 
    -9.413952e-09, -2.784304e-09, 4.168896e-09, 1.132514e-08, -1.482101e-08, 
    2.730495e-08, 1.395483e-09, -1.055616e-08, -2.713989e-08, -2.059414e-08, 
    -8.689995e-09, 7.241533e-08, 1.110777e-08, 1.080866e-08, 3.93984e-08, 
    -1.790568e-10, 1.780472e-08, -3.886998e-08, -1.139927e-08, -1.923968e-08, 
    5.208346e-08, -3.451623e-08, -5.452333e-07, 2.985112e-07, 3.554419e-09, 
    3.153426e-07, -2.364445e-08, 5.942866e-09, -2.173158e-08, 5.566277e-08, 
    -9.284143e-08, 3.360742e-08, -1.155925e-08, -9.014347e-09, -2.156401e-08, 
    -3.428056e-08, 2.278543e-07, 2.947266e-07, -1.621374e-08, -2.590546e-09, 
    9.200639e-08, -1.971864e-08, 1.255903e-08, 3.164669e-08, 4.284343e-08, 
    -6.204175e-09, -4.578874e-08, -6.461836e-09, -1.619182e-08, 
    -1.069934e-08, 1.009073e-08, 8.346319e-09, 1.426861e-08, -3.210114e-07, 
    2.282122e-08, 6.52235e-08, -1.216438e-08, -1.017744e-07, 2.051979e-08, 
    1.255933e-08, -4.61082e-08, -8.120571e-08, -2.279876e-09, 1.615797e-08, 
    3.36132e-08, -4.625804e-09, 4.674341e-08, 6.023981e-10, 2.10127e-10, 
    4.102276e-08, -3.628497e-08, 1.055666e-08, 3.814318e-08, 8.30596e-09, 
    -5.610002e-08, 6.030598e-08, -8.633151e-09, 3.536093e-08, -2.108474e-08, 
    2.193792e-08, -2.885452e-08, 4.869639e-08, 2.749772e-09, -6.162873e-09, 
    1.441754e-08, 5.674932e-08, -3.652224e-08, 3.115747e-08, -2.796696e-08, 
    -1.822537e-09, 2.696277e-08, 4.56727e-08, -8.743768e-08, 4.056915e-09, 
    -1.089295e-07, -2.5796e-08, -9.951623e-08, -3.925845e-08, -8.012648e-10, 
    8.720917e-10, -1.458898e-08, -6.338041e-10, 8.856318e-09, 6.307346e-10, 
    -5.400432e-08, -4.183107e-10, -1.468464e-08, 1.071395e-08, 4.246175e-09, 
    -9.441692e-10 ;
}
