netcdf sos_Omon_exAA03_historical_r3i1p1_185001-200512_box {
dimensions:
	x = 20 ;
	y = 20 ;
	nv4 = 4 ;
	time = UNLIMITED ; // (4 currently)
	bnds = 2 ;
variables:
	float lon(y, x) ;
		lon:standard_name = "longitude" ;
		lon:long_name = "longitude coordinate" ;
		lon:units = "degrees_east" ;
		lon:_CoordinateAxisType = "Lon" ;
		lon:bounds = "lon_bnds" ;
	float lon_bnds(y, x, nv4) ;
	float lat(y, x) ;
		lat:standard_name = "latitude" ;
		lat:long_name = "latitude coordinate" ;
		lat:units = "degrees_north" ;
		lat:_CoordinateAxisType = "Lat" ;
		lat:bounds = "lat_bnds" ;
	float lat_bnds(y, x, nv4) ;
	double time(time) ;
		time:standard_name = "time" ;
		time:long_name = "time" ;
		time:bounds = "time_bnds" ;
		time:units = "days since 1800-1-1 00:00:00" ;
		time:calendar = "365_day" ;
		time:axis = "T" ;
	double time_bnds(time, bnds) ;
	float sos(time, y, x) ;
		sos:standard_name = "sea_surface_salinity" ;
		sos:long_name = "Sea Surface Salinity" ;
		sos:units = "psu" ;
		sos:coordinates = "lat lon" ;
		sos:_FillValue = 1.e+20f ;
		sos:missing_value = 1.e+20f ;
		sos:original_name = "sss" ;
		sos:cell_methods = "time: mean" ;
		sos:history = "2011-07-16T20:41:19Z altered by CMOR: replaced missing value flag (1e+20) with standard missing value (1e+20). 2011-07-16T20:41:19Z altered by CMOR: Converted type from \'d\' to \'f\'." ;
		sos:associated_files = "baseURL: http://cmip-pcmdi.llnl.gov/CMIP5/dataLocation gridspecFile: gridspec_ocean_fx_NorESM1-M_historical_r0i0p0.nc areacello: areacello_fx_NorESM1-M_historical_r0i0p0.nc" ;

// global attributes:
		:CDI = "Climate Data Interface version ?? (http://mpimet.mpg.de/cdi)" ;
		:Conventions = "CF-1.4" ;
		:history = "reset by cdo to create anonymous sample file" ;
		:source = "201707_compliance_checker_evaluation/work/p1.py" ;
		:institution = "CEDA" ;
		:institute_id = "CEDA" ;
		:experiment_id = "historical" ;
		:model_id = "exAA03" ;
		:forcing = "GHG, SA, Oz, Sl, Vl, BC, OC" ;
		:parent_experiment_id = "piControl" ;
		:parent_experiment_rip = "r1i1p1" ;
		:branch_time = 277035. ;
		:contact = "none" ;
		:initialization_method = 1 ;
		:physics_version = 1 ;
		:tracking_id = "47bb552c-cb54-4d85-9fb8-fc524fa2ae21" ;
		:product = "output" ;
		:experiment = "historical" ;
		:frequency = "mon" ;
		:creation_date = "2011-07-16T20:41:19Z" ;
		:project_id = "CMIP5" ;
		:table_id = "Table Omon (27 April 2011) 340eddd4fd838d90fa9ffe1345ecbd73" ;
		:title = "Dummy file with known metadata errors" ;
		:parent_experiment = "pre-industrial control" ;
		:modeling_realm = "ocean" ;
		:realization = 3 ;
		:cmor_version = "2.7.1" ;
		:comment = "this is a sample file with known metadata errors" ;
		:CDO = "Climate Data Operators version 1.7.0 (http://mpimet.mpg.de/cdo)" ;
data:

 lon =
  320.5625, 321.6875, 322.8125, 323.9375, 325.0625, 326.1875, 327.3125, 
    328.4375, 329.5625, 330.6875, 331.8125, 332.9375, 334.0625, 335.1875, 
    336.3125, 337.4375, 338.5625, 339.6875, 340.8125, 341.9375,
  320.5625, 321.6875, 322.8125, 323.9375, 325.0625, 326.1875, 327.3125, 
    328.4375, 329.5625, 330.6875, 331.8125, 332.9375, 334.0625, 335.1875, 
    336.3125, 337.4375, 338.5625, 339.6875, 340.8125, 341.9375,
  320.5625, 321.6875, 322.8125, 323.9375, 325.0625, 326.1875, 327.3125, 
    328.4375, 329.5625, 330.6875, 331.8125, 332.9375, 334.0625, 335.1875, 
    336.3125, 337.4375, 338.5625, 339.6875, 340.8125, 341.9375,
  320.5625, 321.6875, 322.8125, 323.9375, 325.0625, 326.1875, 327.3125, 
    328.4375, 329.5625, 330.6875, 331.8125, 332.9375, 334.0625, 335.1875, 
    336.3125, 337.4375, 338.5625, 339.6875, 340.8125, 341.9375,
  320.5625, 321.6875, 322.8125, 323.9375, 325.0625, 326.1875, 327.3125, 
    328.4375, 329.5625, 330.6875, 331.8125, 332.9375, 334.0625, 335.1875, 
    336.3125, 337.4375, 338.5625, 339.6875, 340.8125, 341.9375,
  320.5625, 321.6875, 322.8125, 323.9375, 325.0625, 326.1875, 327.3125, 
    328.4375, 329.5625, 330.6875, 331.8125, 332.9375, 334.0625, 335.1875, 
    336.3125, 337.4375, 338.5625, 339.6875, 340.8125, 341.9375,
  320.5625, 321.6875, 322.8125, 323.9375, 325.0625, 326.1875, 327.3125, 
    328.4375, 329.5625, 330.6875, 331.8125, 332.9375, 334.0625, 335.1875, 
    336.3125, 337.4375, 338.5625, 339.6875, 340.8125, 341.9375,
  320.5625, 321.6875, 322.8125, 323.9375, 325.0625, 326.1875, 327.3125, 
    328.4375, 329.5625, 330.6875, 331.8125, 332.9375, 334.0625, 335.1875, 
    336.3125, 337.4375, 338.5625, 339.6875, 340.8125, 341.9375,
  320.5625, 321.6875, 322.8125, 323.9375, 325.0625, 326.1875, 327.3125, 
    328.4375, 329.5625, 330.6875, 331.8125, 332.9375, 334.0625, 335.1875, 
    336.3125, 337.4375, 338.5625, 339.6875, 340.8125, 341.9375,
  320.5625, 321.6875, 322.8125, 323.9375, 325.0625, 326.1875, 327.3125, 
    328.4375, 329.5625, 330.6875, 331.8125, 332.9375, 334.0625, 335.1875, 
    336.3125, 337.4375, 338.5625, 339.6875, 340.8125, 341.9375,
  320.5625, 321.6875, 322.8125, 323.9375, 325.0625, 326.1875, 327.3125, 
    328.4375, 329.5625, 330.6875, 331.8125, 332.9375, 334.0625, 335.1875, 
    336.3125, 337.4375, 338.5625, 339.6875, 340.8125, 341.9375,
  320.5625, 321.6875, 322.8125, 323.9375, 325.0625, 326.1875, 327.3125, 
    328.4375, 329.5625, 330.6875, 331.8125, 332.9375, 334.0625, 335.1875, 
    336.3125, 337.4375, 338.5625, 339.6875, 340.8125, 341.9375,
  320.5625, 321.6875, 322.8125, 323.9375, 325.0625, 326.1875, 327.3125, 
    328.4375, 329.5625, 330.6875, 331.8125, 332.9375, 334.0625, 335.1875, 
    336.3125, 337.4375, 338.5625, 339.6875, 340.8125, 341.9375,
  320.5625, 321.6875, 322.8125, 323.9375, 325.0625, 326.1875, 327.3125, 
    328.4375, 329.5625, 330.6875, 331.8125, 332.9375, 334.0625, 335.1875, 
    336.3125, 337.4375, 338.5625, 339.6875, 340.8125, 341.9375,
  320.5625, 321.6875, 322.8125, 323.9375, 325.0625, 326.1875, 327.3125, 
    328.4375, 329.5625, 330.6875, 331.8125, 332.9375, 334.0625, 335.1875, 
    336.3125, 337.4375, 338.5625, 339.6875, 340.8125, 341.9375,
  320.5625, 321.6875, 322.8125, 323.9375, 325.0625, 326.1875, 327.3125, 
    328.4375, 329.5625, 330.6875, 331.8125, 332.9375, 334.0625, 335.1875, 
    336.3125, 337.4375, 338.5625, 339.6875, 340.8125, 341.9375,
  320.5625, 321.6875, 322.8125, 323.9375, 325.0625, 326.1875, 327.3125, 
    328.4375, 329.5625, 330.6875, 331.8125, 332.9375, 334.0625, 335.1875, 
    336.3125, 337.4375, 338.5625, 339.6875, 340.8125, 341.9375,
  320.5625, 321.6875, 322.8125, 323.9375, 325.0625, 326.1875, 327.3125, 
    328.4375, 329.5625, 330.6875, 331.8125, 332.9375, 334.0625, 335.1875, 
    336.3125, 337.4375, 338.5625, 339.6875, 340.8125, 341.9375,
  320.5625, 321.6875, 322.8125, 323.9375, 325.0625, 326.1875, 327.3125, 
    328.4375, 329.5625, 330.6875, 331.8125, 332.9375, 334.0625, 335.1875, 
    336.3125, 337.4375, 338.5625, 339.6875, 340.8125, 341.9375,
  320.5625, 321.6875, 322.8125, 323.9375, 325.0625, 326.1875, 327.3125, 
    328.4375, 329.5625, 330.6875, 331.8125, 332.9375, 334.0625, 335.1875, 
    336.3125, 337.4375, 338.5625, 339.6875, 340.8125, 341.9375 ;

 lon_bnds =
  320, 321.125, 321.125, 320,
  321.125, 322.25, 322.25, 321.125,
  322.25, 323.375, 323.375, 322.25,
  323.375, 324.5, 324.5, 323.375,
  324.5, 325.625, 325.625, 324.5,
  325.625, 326.75, 326.75, 325.625,
  326.75, 327.875, 327.875, 326.75,
  327.875, 329, 329, 327.875,
  329, 330.125, 330.125, 329,
  330.125, 331.25, 331.25, 330.125,
  331.25, 332.375, 332.375, 331.25,
  332.375, 333.5, 333.5, 332.375,
  333.5, 334.625, 334.625, 333.5,
  334.625, 335.75, 335.75, 334.625,
  335.75, 336.875, 336.875, 335.75,
  336.875, 338, 338, 336.875,
  338, 339.125, 339.125, 338,
  339.125, 340.25, 340.25, 339.125,
  340.25, 341.375, 341.375, 340.25,
  341.375, 342.5, 342.5, 341.375,
  320, 321.125, 321.125, 320,
  321.125, 322.25, 322.25, 321.125,
  322.25, 323.375, 323.375, 322.25,
  323.375, 324.5, 324.5, 323.375,
  324.5, 325.625, 325.625, 324.5,
  325.625, 326.75, 326.75, 325.625,
  326.75, 327.875, 327.875, 326.75,
  327.875, 329, 329, 327.875,
  329, 330.125, 330.125, 329,
  330.125, 331.25, 331.25, 330.125,
  331.25, 332.375, 332.375, 331.25,
  332.375, 333.5, 333.5, 332.375,
  333.5, 334.625, 334.625, 333.5,
  334.625, 335.75, 335.75, 334.625,
  335.75, 336.875, 336.875, 335.75,
  336.875, 338, 338, 336.875,
  338, 339.125, 339.125, 338,
  339.125, 340.25, 340.25, 339.125,
  340.25, 341.375, 341.375, 340.25,
  341.375, 342.5, 342.5, 341.375,
  320, 321.125, 321.125, 320,
  321.125, 322.25, 322.25, 321.125,
  322.25, 323.375, 323.375, 322.25,
  323.375, 324.5, 324.5, 323.375,
  324.5, 325.625, 325.625, 324.5,
  325.625, 326.75, 326.75, 325.625,
  326.75, 327.875, 327.875, 326.75,
  327.875, 329, 329, 327.875,
  329, 330.125, 330.125, 329,
  330.125, 331.25, 331.25, 330.125,
  331.25, 332.375, 332.375, 331.25,
  332.375, 333.5, 333.5, 332.375,
  333.5, 334.625, 334.625, 333.5,
  334.625, 335.75, 335.75, 334.625,
  335.75, 336.875, 336.875, 335.75,
  336.875, 338, 338, 336.875,
  338, 339.125, 339.125, 338,
  339.125, 340.25, 340.25, 339.125,
  340.25, 341.375, 341.375, 340.25,
  341.375, 342.5, 342.5, 341.375,
  320, 321.125, 321.125, 320,
  321.125, 322.25, 322.25, 321.125,
  322.25, 323.375, 323.375, 322.25,
  323.375, 324.5, 324.5, 323.375,
  324.5, 325.625, 325.625, 324.5,
  325.625, 326.75, 326.75, 325.625,
  326.75, 327.875, 327.875, 326.75,
  327.875, 329, 329, 327.875,
  329, 330.125, 330.125, 329,
  330.125, 331.25, 331.25, 330.125,
  331.25, 332.375, 332.375, 331.25,
  332.375, 333.5, 333.5, 332.375,
  333.5, 334.625, 334.625, 333.5,
  334.625, 335.75, 335.75, 334.625,
  335.75, 336.875, 336.875, 335.75,
  336.875, 338, 338, 336.875,
  338, 339.125, 339.125, 338,
  339.125, 340.25, 340.25, 339.125,
  340.25, 341.375, 341.375, 340.25,
  341.375, 342.5, 342.5, 341.375,
  320, 321.125, 321.125, 320,
  321.125, 322.25, 322.25, 321.125,
  322.25, 323.375, 323.375, 322.25,
  323.375, 324.5, 324.5, 323.375,
  324.5, 325.625, 325.625, 324.5,
  325.625, 326.75, 326.75, 325.625,
  326.75, 327.875, 327.875, 326.75,
  327.875, 329, 329, 327.875,
  329, 330.125, 330.125, 329,
  330.125, 331.25, 331.25, 330.125,
  331.25, 332.375, 332.375, 331.25,
  332.375, 333.5, 333.5, 332.375,
  333.5, 334.625, 334.625, 333.5,
  334.625, 335.75, 335.75, 334.625,
  335.75, 336.875, 336.875, 335.75,
  336.875, 338, 338, 336.875,
  338, 339.125, 339.125, 338,
  339.125, 340.25, 340.25, 339.125,
  340.25, 341.375, 341.375, 340.25,
  341.375, 342.5, 342.5, 341.375,
  320, 321.125, 321.125, 320,
  321.125, 322.25, 322.25, 321.125,
  322.25, 323.375, 323.375, 322.25,
  323.375, 324.5, 324.5, 323.375,
  324.5, 325.625, 325.625, 324.5,
  325.625, 326.75, 326.75, 325.625,
  326.75, 327.875, 327.875, 326.75,
  327.875, 329, 329, 327.875,
  329, 330.125, 330.125, 329,
  330.125, 331.25, 331.25, 330.125,
  331.25, 332.375, 332.375, 331.25,
  332.375, 333.5, 333.5, 332.375,
  333.5, 334.625, 334.625, 333.5,
  334.625, 335.75, 335.75, 334.625,
  335.75, 336.875, 336.875, 335.75,
  336.875, 338, 338, 336.875,
  338, 339.125, 339.125, 338,
  339.125, 340.25, 340.25, 339.125,
  340.25, 341.375, 341.375, 340.25,
  341.375, 342.5, 342.5, 341.375,
  320, 321.125, 321.125, 320,
  321.125, 322.25, 322.25, 321.125,
  322.25, 323.375, 323.375, 322.25,
  323.375, 324.5, 324.5, 323.375,
  324.5, 325.625, 325.625, 324.5,
  325.625, 326.75, 326.75, 325.625,
  326.75, 327.875, 327.875, 326.75,
  327.875, 329, 329, 327.875,
  329, 330.125, 330.125, 329,
  330.125, 331.25, 331.25, 330.125,
  331.25, 332.375, 332.375, 331.25,
  332.375, 333.5, 333.5, 332.375,
  333.5, 334.625, 334.625, 333.5,
  334.625, 335.75, 335.75, 334.625,
  335.75, 336.875, 336.875, 335.75,
  336.875, 338, 338, 336.875,
  338, 339.125, 339.125, 338,
  339.125, 340.25, 340.25, 339.125,
  340.25, 341.375, 341.375, 340.25,
  341.375, 342.5, 342.5, 341.375,
  320, 321.125, 321.125, 320,
  321.125, 322.25, 322.25, 321.125,
  322.25, 323.375, 323.375, 322.25,
  323.375, 324.5, 324.5, 323.375,
  324.5, 325.625, 325.625, 324.5,
  325.625, 326.75, 326.75, 325.625,
  326.75, 327.875, 327.875, 326.75,
  327.875, 329, 329, 327.875,
  329, 330.125, 330.125, 329,
  330.125, 331.25, 331.25, 330.125,
  331.25, 332.375, 332.375, 331.25,
  332.375, 333.5, 333.5, 332.375,
  333.5, 334.625, 334.625, 333.5,
  334.625, 335.75, 335.75, 334.625,
  335.75, 336.875, 336.875, 335.75,
  336.875, 338, 338, 336.875,
  338, 339.125, 339.125, 338,
  339.125, 340.25, 340.25, 339.125,
  340.25, 341.375, 341.375, 340.25,
  341.375, 342.5, 342.5, 341.375,
  320, 321.125, 321.125, 320,
  321.125, 322.25, 322.25, 321.125,
  322.25, 323.375, 323.375, 322.25,
  323.375, 324.5, 324.5, 323.375,
  324.5, 325.625, 325.625, 324.5,
  325.625, 326.75, 326.75, 325.625,
  326.75, 327.875, 327.875, 326.75,
  327.875, 329, 329, 327.875,
  329, 330.125, 330.125, 329,
  330.125, 331.25, 331.25, 330.125,
  331.25, 332.375, 332.375, 331.25,
  332.375, 333.5, 333.5, 332.375,
  333.5, 334.625, 334.625, 333.5,
  334.625, 335.75, 335.75, 334.625,
  335.75, 336.875, 336.875, 335.75,
  336.875, 338, 338, 336.875,
  338, 339.125, 339.125, 338,
  339.125, 340.25, 340.25, 339.125,
  340.25, 341.375, 341.375, 340.25,
  341.375, 342.5, 342.5, 341.375,
  320, 321.125, 321.125, 320,
  321.125, 322.25, 322.25, 321.125,
  322.25, 323.375, 323.375, 322.25,
  323.375, 324.5, 324.5, 323.375,
  324.5, 325.625, 325.625, 324.5,
  325.625, 326.75, 326.75, 325.625,
  326.75, 327.875, 327.875, 326.75,
  327.875, 329, 329, 327.875,
  329, 330.125, 330.125, 329,
  330.125, 331.25, 331.25, 330.125,
  331.25, 332.375, 332.375, 331.25,
  332.375, 333.5, 333.5, 332.375,
  333.5, 334.625, 334.625, 333.5,
  334.625, 335.75, 335.75, 334.625,
  335.75, 336.875, 336.875, 335.75,
  336.875, 338, 338, 336.875,
  338, 339.125, 339.125, 338,
  339.125, 340.25, 340.25, 339.125,
  340.25, 341.375, 341.375, 340.25,
  341.375, 342.5, 342.5, 341.375,
  320, 321.125, 321.125, 320,
  321.125, 322.25, 322.25, 321.125,
  322.25, 323.375, 323.375, 322.25,
  323.375, 324.5, 324.5, 323.375,
  324.5, 325.625, 325.625, 324.5,
  325.625, 326.75, 326.75, 325.625,
  326.75, 327.875, 327.875, 326.75,
  327.875, 329, 329, 327.875,
  329, 330.125, 330.125, 329,
  330.125, 331.25, 331.25, 330.125,
  331.25, 332.375, 332.375, 331.25,
  332.375, 333.5, 333.5, 332.375,
  333.5, 334.625, 334.625, 333.5,
  334.625, 335.75, 335.75, 334.625,
  335.75, 336.875, 336.875, 335.75,
  336.875, 338, 338, 336.875,
  338, 339.125, 339.125, 338,
  339.125, 340.25, 340.25, 339.125,
  340.25, 341.375, 341.375, 340.25,
  341.375, 342.5, 342.5, 341.375,
  320, 321.125, 321.125, 320,
  321.125, 322.25, 322.25, 321.125,
  322.25, 323.375, 323.375, 322.25,
  323.375, 324.5, 324.5, 323.375,
  324.5, 325.625, 325.625, 324.5,
  325.625, 326.75, 326.75, 325.625,
  326.75, 327.875, 327.875, 326.75,
  327.875, 329, 329, 327.875,
  329, 330.125, 330.125, 329,
  330.125, 331.25, 331.25, 330.125,
  331.25, 332.375, 332.375, 331.25,
  332.375, 333.5, 333.5, 332.375,
  333.5, 334.625, 334.625, 333.5,
  334.625, 335.75, 335.75, 334.625,
  335.75, 336.875, 336.875, 335.75,
  336.875, 338, 338, 336.875,
  338, 339.125, 339.125, 338,
  339.125, 340.25, 340.25, 339.125,
  340.25, 341.375, 341.375, 340.25,
  341.375, 342.5, 342.5, 341.375,
  320, 321.125, 321.125, 320,
  321.125, 322.25, 322.25, 321.125,
  322.25, 323.375, 323.375, 322.25,
  323.375, 324.5, 324.5, 323.375,
  324.5, 325.625, 325.625, 324.5,
  325.625, 326.75, 326.75, 325.625,
  326.75, 327.875, 327.875, 326.75,
  327.875, 329, 329, 327.875,
  329, 330.125, 330.125, 329,
  330.125, 331.25, 331.25, 330.125,
  331.25, 332.375, 332.375, 331.25,
  332.375, 333.5, 333.5, 332.375,
  333.5, 334.625, 334.625, 333.5,
  334.625, 335.75, 335.75, 334.625,
  335.75, 336.875, 336.875, 335.75,
  336.875, 338, 338, 336.875,
  338, 339.125, 339.125, 338,
  339.125, 340.25, 340.25, 339.125,
  340.25, 341.375, 341.375, 340.25,
  341.375, 342.5, 342.5, 341.375,
  320, 321.125, 321.125, 320,
  321.125, 322.25, 322.25, 321.125,
  322.25, 323.375, 323.375, 322.25,
  323.375, 324.5, 324.5, 323.375,
  324.5, 325.625, 325.625, 324.5,
  325.625, 326.75, 326.75, 325.625,
  326.75, 327.875, 327.875, 326.75,
  327.875, 329, 329, 327.875,
  329, 330.125, 330.125, 329,
  330.125, 331.25, 331.25, 330.125,
  331.25, 332.375, 332.375, 331.25,
  332.375, 333.5, 333.5, 332.375,
  333.5, 334.625, 334.625, 333.5,
  334.625, 335.75, 335.75, 334.625,
  335.75, 336.875, 336.875, 335.75,
  336.875, 338, 338, 336.875,
  338, 339.125, 339.125, 338,
  339.125, 340.25, 340.25, 339.125,
  340.25, 341.375, 341.375, 340.25,
  341.375, 342.5, 342.5, 341.375,
  320, 321.125, 321.125, 320,
  321.125, 322.25, 322.25, 321.125,
  322.25, 323.375, 323.375, 322.25,
  323.375, 324.5, 324.5, 323.375,
  324.5, 325.625, 325.625, 324.5,
  325.625, 326.75, 326.75, 325.625,
  326.75, 327.875, 327.875, 326.75,
  327.875, 329, 329, 327.875,
  329, 330.125, 330.125, 329,
  330.125, 331.25, 331.25, 330.125,
  331.25, 332.375, 332.375, 331.25,
  332.375, 333.5, 333.5, 332.375,
  333.5, 334.625, 334.625, 333.5,
  334.625, 335.75, 335.75, 334.625,
  335.75, 336.875, 336.875, 335.75,
  336.875, 338, 338, 336.875,
  338, 339.125, 339.125, 338,
  339.125, 340.25, 340.25, 339.125,
  340.25, 341.375, 341.375, 340.25,
  341.375, 342.5, 342.5, 341.375,
  320, 321.125, 321.125, 320,
  321.125, 322.25, 322.25, 321.125,
  322.25, 323.375, 323.375, 322.25,
  323.375, 324.5, 324.5, 323.375,
  324.5, 325.625, 325.625, 324.5,
  325.625, 326.75, 326.75, 325.625,
  326.75, 327.875, 327.875, 326.75,
  327.875, 329, 329, 327.875,
  329, 330.125, 330.125, 329,
  330.125, 331.25, 331.25, 330.125,
  331.25, 332.375, 332.375, 331.25,
  332.375, 333.5, 333.5, 332.375,
  333.5, 334.625, 334.625, 333.5,
  334.625, 335.75, 335.75, 334.625,
  335.75, 336.875, 336.875, 335.75,
  336.875, 338, 338, 336.875,
  338, 339.125, 339.125, 338,
  339.125, 340.25, 340.25, 339.125,
  340.25, 341.375, 341.375, 340.25,
  341.375, 342.5, 342.5, 341.375,
  320, 321.125, 321.125, 320,
  321.125, 322.25, 322.25, 321.125,
  322.25, 323.375, 323.375, 322.25,
  323.375, 324.5, 324.5, 323.375,
  324.5, 325.625, 325.625, 324.5,
  325.625, 326.75, 326.75, 325.625,
  326.75, 327.875, 327.875, 326.75,
  327.875, 329, 329, 327.875,
  329, 330.125, 330.125, 329,
  330.125, 331.25, 331.25, 330.125,
  331.25, 332.375, 332.375, 331.25,
  332.375, 333.5, 333.5, 332.375,
  333.5, 334.625, 334.625, 333.5,
  334.625, 335.75, 335.75, 334.625,
  335.75, 336.875, 336.875, 335.75,
  336.875, 338, 338, 336.875,
  338, 339.125, 339.125, 338,
  339.125, 340.25, 340.25, 339.125,
  340.25, 341.375, 341.375, 340.25,
  341.375, 342.5, 342.5, 341.375,
  320, 321.125, 321.125, 320,
  321.125, 322.25, 322.25, 321.125,
  322.25, 323.375, 323.375, 322.25,
  323.375, 324.5, 324.5, 323.375,
  324.5, 325.625, 325.625, 324.5,
  325.625, 326.75, 326.75, 325.625,
  326.75, 327.875, 327.875, 326.75,
  327.875, 329, 329, 327.875,
  329, 330.125, 330.125, 329,
  330.125, 331.25, 331.25, 330.125,
  331.25, 332.375, 332.375, 331.25,
  332.375, 333.5, 333.5, 332.375,
  333.5, 334.625, 334.625, 333.5,
  334.625, 335.75, 335.75, 334.625,
  335.75, 336.875, 336.875, 335.75,
  336.875, 338, 338, 336.875,
  338, 339.125, 339.125, 338,
  339.125, 340.25, 340.25, 339.125,
  340.25, 341.375, 341.375, 340.25,
  341.375, 342.5, 342.5, 341.375,
  320, 321.125, 321.125, 320,
  321.125, 322.25, 322.25, 321.125,
  322.25, 323.375, 323.375, 322.25,
  323.375, 324.5, 324.5, 323.375,
  324.5, 325.625, 325.625, 324.5,
  325.625, 326.75, 326.75, 325.625,
  326.75, 327.875, 327.875, 326.75,
  327.875, 329, 329, 327.875,
  329, 330.125, 330.125, 329,
  330.125, 331.25, 331.25, 330.125,
  331.25, 332.375, 332.375, 331.25,
  332.375, 333.5, 333.5, 332.375,
  333.5, 334.625, 334.625, 333.5,
  334.625, 335.75, 335.75, 334.625,
  335.75, 336.875, 336.875, 335.75,
  336.875, 338, 338, 336.875,
  338, 339.125, 339.125, 338,
  339.125, 340.25, 340.25, 339.125,
  340.25, 341.375, 341.375, 340.25,
  341.375, 342.5, 342.5, 341.375,
  320, 321.125, 321.125, 320,
  321.125, 322.25, 322.25, 321.125,
  322.25, 323.375, 323.375, 322.25,
  323.375, 324.5, 324.5, 323.375,
  324.5, 325.625, 325.625, 324.5,
  325.625, 326.75, 326.75, 325.625,
  326.75, 327.875, 327.875, 326.75,
  327.875, 329, 329, 327.875,
  329, 330.125, 330.125, 329,
  330.125, 331.25, 331.25, 330.125,
  331.25, 332.375, 332.375, 331.25,
  332.375, 333.5, 333.5, 332.375,
  333.5, 334.625, 334.625, 333.5,
  334.625, 335.75, 335.75, 334.625,
  335.75, 336.875, 336.875, 335.75,
  336.875, 338, 338, 336.875,
  338, 339.125, 339.125, 338,
  339.125, 340.25, 340.25, 339.125,
  340.25, 341.375, 341.375, 340.25,
  341.375, 342.5, 342.5, 341.375 ;

 lat =
  -79.22052, -79.22052, -79.22052, -79.22052, -79.22052, -79.22052, 
    -79.22052, -79.22052, -79.22052, -79.22052, -79.22052, -79.22052, 
    -79.22052, -79.22052, -79.22052, -79.22052, -79.22052, -79.22052, 
    -79.22052, -79.22052,
  -78.68631, -78.68631, -78.68631, -78.68631, -78.68631, -78.68631, 
    -78.68631, -78.68631, -78.68631, -78.68631, -78.68631, -78.68631, 
    -78.68631, -78.68631, -78.68631, -78.68631, -78.68631, -78.68631, 
    -78.68631, -78.68631,
  -78.15209, -78.15209, -78.15209, -78.15209, -78.15209, -78.15209, 
    -78.15209, -78.15209, -78.15209, -78.15209, -78.15209, -78.15209, 
    -78.15209, -78.15209, -78.15209, -78.15209, -78.15209, -78.15209, 
    -78.15209, -78.15209,
  -77.61787, -77.61787, -77.61787, -77.61787, -77.61787, -77.61787, 
    -77.61787, -77.61787, -77.61787, -77.61787, -77.61787, -77.61787, 
    -77.61787, -77.61787, -77.61787, -77.61787, -77.61787, -77.61787, 
    -77.61787, -77.61787,
  -77.08366, -77.08366, -77.08366, -77.08366, -77.08366, -77.08366, 
    -77.08366, -77.08366, -77.08366, -77.08366, -77.08366, -77.08366, 
    -77.08366, -77.08366, -77.08366, -77.08366, -77.08366, -77.08366, 
    -77.08366, -77.08366,
  -76.54944, -76.54944, -76.54944, -76.54944, -76.54944, -76.54944, 
    -76.54944, -76.54944, -76.54944, -76.54944, -76.54944, -76.54944, 
    -76.54944, -76.54944, -76.54944, -76.54944, -76.54944, -76.54944, 
    -76.54944, -76.54944,
  -76.01522, -76.01522, -76.01522, -76.01522, -76.01522, -76.01522, 
    -76.01522, -76.01522, -76.01522, -76.01522, -76.01522, -76.01522, 
    -76.01522, -76.01522, -76.01522, -76.01522, -76.01522, -76.01522, 
    -76.01522, -76.01522,
  -75.481, -75.481, -75.481, -75.481, -75.481, -75.481, -75.481, -75.481, 
    -75.481, -75.481, -75.481, -75.481, -75.481, -75.481, -75.481, -75.481, 
    -75.481, -75.481, -75.481, -75.481,
  -74.94678, -74.94678, -74.94678, -74.94678, -74.94678, -74.94678, 
    -74.94678, -74.94678, -74.94678, -74.94678, -74.94678, -74.94678, 
    -74.94678, -74.94678, -74.94678, -74.94678, -74.94678, -74.94678, 
    -74.94678, -74.94678,
  -74.41257, -74.41257, -74.41257, -74.41257, -74.41257, -74.41257, 
    -74.41257, -74.41257, -74.41257, -74.41257, -74.41257, -74.41257, 
    -74.41257, -74.41257, -74.41257, -74.41257, -74.41257, -74.41257, 
    -74.41257, -74.41257,
  -73.87835, -73.87835, -73.87835, -73.87835, -73.87835, -73.87835, 
    -73.87835, -73.87835, -73.87835, -73.87835, -73.87835, -73.87835, 
    -73.87835, -73.87835, -73.87835, -73.87835, -73.87835, -73.87835, 
    -73.87835, -73.87835,
  -73.34413, -73.34413, -73.34413, -73.34413, -73.34413, -73.34413, 
    -73.34413, -73.34413, -73.34413, -73.34413, -73.34413, -73.34413, 
    -73.34413, -73.34413, -73.34413, -73.34413, -73.34413, -73.34413, 
    -73.34413, -73.34413,
  -72.80991, -72.80991, -72.80991, -72.80991, -72.80991, -72.80991, 
    -72.80991, -72.80991, -72.80991, -72.80991, -72.80991, -72.80991, 
    -72.80991, -72.80991, -72.80991, -72.80991, -72.80991, -72.80991, 
    -72.80991, -72.80991,
  -72.2757, -72.2757, -72.2757, -72.2757, -72.2757, -72.2757, -72.2757, 
    -72.2757, -72.2757, -72.2757, -72.2757, -72.2757, -72.2757, -72.2757, 
    -72.2757, -72.2757, -72.2757, -72.2757, -72.2757, -72.2757,
  -71.74148, -71.74148, -71.74148, -71.74148, -71.74148, -71.74148, 
    -71.74148, -71.74148, -71.74148, -71.74148, -71.74148, -71.74148, 
    -71.74148, -71.74148, -71.74148, -71.74148, -71.74148, -71.74148, 
    -71.74148, -71.74148,
  -71.20726, -71.20726, -71.20726, -71.20726, -71.20726, -71.20726, 
    -71.20726, -71.20726, -71.20726, -71.20726, -71.20726, -71.20726, 
    -71.20726, -71.20726, -71.20726, -71.20726, -71.20726, -71.20726, 
    -71.20726, -71.20726,
  -70.67303, -70.67303, -70.67303, -70.67303, -70.67303, -70.67303, 
    -70.67303, -70.67303, -70.67303, -70.67303, -70.67303, -70.67303, 
    -70.67303, -70.67303, -70.67303, -70.67303, -70.67303, -70.67303, 
    -70.67303, -70.67303,
  -70.13882, -70.13882, -70.13882, -70.13882, -70.13882, -70.13882, 
    -70.13882, -70.13882, -70.13882, -70.13882, -70.13882, -70.13882, 
    -70.13882, -70.13882, -70.13882, -70.13882, -70.13882, -70.13882, 
    -70.13882, -70.13882,
  -69.6046, -69.6046, -69.6046, -69.6046, -69.6046, -69.6046, -69.6046, 
    -69.6046, -69.6046, -69.6046, -69.6046, -69.6046, -69.6046, -69.6046, 
    -69.6046, -69.6046, -69.6046, -69.6046, -69.6046, -69.6046,
  -69.07037, -69.07037, -69.07037, -69.07037, -69.07037, -69.07037, 
    -69.07037, -69.07037, -69.07037, -69.07037, -69.07037, -69.07037, 
    -69.07037, -69.07037, -69.07037, -69.07037, -69.07037, -69.07037, 
    -69.07037, -69.07037 ;

 lat_bnds =
  -79.48714, -79.48714, -78.9529, -78.9529,
  -79.48714, -79.48714, -78.9529, -78.9529,
  -79.48714, -79.48714, -78.9529, -78.9529,
  -79.48714, -79.48714, -78.9529, -78.9529,
  -79.48714, -79.48714, -78.9529, -78.9529,
  -79.48714, -79.48714, -78.9529, -78.9529,
  -79.48714, -79.48714, -78.9529, -78.9529,
  -79.48714, -79.48714, -78.9529, -78.9529,
  -79.48714, -79.48714, -78.9529, -78.9529,
  -79.48714, -79.48714, -78.9529, -78.9529,
  -79.48714, -79.48714, -78.9529, -78.9529,
  -79.48714, -79.48714, -78.9529, -78.9529,
  -79.48714, -79.48714, -78.9529, -78.9529,
  -79.48714, -79.48714, -78.9529, -78.9529,
  -79.48714, -79.48714, -78.9529, -78.9529,
  -79.48714, -79.48714, -78.9529, -78.9529,
  -79.48714, -79.48714, -78.9529, -78.9529,
  -79.48714, -79.48714, -78.9529, -78.9529,
  -79.48714, -79.48714, -78.9529, -78.9529,
  -79.48714, -79.48714, -78.9529, -78.9529,
  -78.9529, -78.9529, -78.41866, -78.41866,
  -78.9529, -78.9529, -78.41866, -78.41866,
  -78.9529, -78.9529, -78.41866, -78.41866,
  -78.9529, -78.9529, -78.41866, -78.41866,
  -78.9529, -78.9529, -78.41866, -78.41866,
  -78.9529, -78.9529, -78.41866, -78.41866,
  -78.9529, -78.9529, -78.41866, -78.41866,
  -78.9529, -78.9529, -78.41866, -78.41866,
  -78.9529, -78.9529, -78.41866, -78.41866,
  -78.9529, -78.9529, -78.41866, -78.41866,
  -78.9529, -78.9529, -78.41866, -78.41866,
  -78.9529, -78.9529, -78.41866, -78.41866,
  -78.9529, -78.9529, -78.41866, -78.41866,
  -78.9529, -78.9529, -78.41866, -78.41866,
  -78.9529, -78.9529, -78.41866, -78.41866,
  -78.9529, -78.9529, -78.41866, -78.41866,
  -78.9529, -78.9529, -78.41866, -78.41866,
  -78.9529, -78.9529, -78.41866, -78.41866,
  -78.9529, -78.9529, -78.41866, -78.41866,
  -78.9529, -78.9529, -78.41866, -78.41866,
  -78.41866, -78.41866, -77.88441, -77.88441,
  -78.41866, -78.41866, -77.88441, -77.88441,
  -78.41866, -78.41866, -77.88441, -77.88441,
  -78.41866, -78.41866, -77.88441, -77.88441,
  -78.41866, -78.41866, -77.88441, -77.88441,
  -78.41866, -78.41866, -77.88441, -77.88441,
  -78.41866, -78.41866, -77.88441, -77.88441,
  -78.41866, -78.41866, -77.88441, -77.88441,
  -78.41866, -78.41866, -77.88441, -77.88441,
  -78.41866, -78.41866, -77.88441, -77.88441,
  -78.41866, -78.41866, -77.88441, -77.88441,
  -78.41866, -78.41866, -77.88441, -77.88441,
  -78.41866, -78.41866, -77.88441, -77.88441,
  -78.41866, -78.41866, -77.88441, -77.88441,
  -78.41866, -78.41866, -77.88441, -77.88441,
  -78.41866, -78.41866, -77.88441, -77.88441,
  -78.41866, -78.41866, -77.88441, -77.88441,
  -78.41866, -78.41866, -77.88441, -77.88441,
  -78.41866, -78.41866, -77.88441, -77.88441,
  -78.41866, -78.41866, -77.88441, -77.88441,
  -77.88441, -77.88441, -77.35017, -77.35017,
  -77.88441, -77.88441, -77.35017, -77.35017,
  -77.88441, -77.88441, -77.35017, -77.35017,
  -77.88441, -77.88441, -77.35017, -77.35017,
  -77.88441, -77.88441, -77.35017, -77.35017,
  -77.88441, -77.88441, -77.35017, -77.35017,
  -77.88441, -77.88441, -77.35017, -77.35017,
  -77.88441, -77.88441, -77.35017, -77.35017,
  -77.88441, -77.88441, -77.35017, -77.35017,
  -77.88441, -77.88441, -77.35017, -77.35017,
  -77.88441, -77.88441, -77.35017, -77.35017,
  -77.88441, -77.88441, -77.35017, -77.35017,
  -77.88441, -77.88441, -77.35017, -77.35017,
  -77.88441, -77.88441, -77.35017, -77.35017,
  -77.88441, -77.88441, -77.35017, -77.35017,
  -77.88441, -77.88441, -77.35017, -77.35017,
  -77.88441, -77.88441, -77.35017, -77.35017,
  -77.88441, -77.88441, -77.35017, -77.35017,
  -77.88441, -77.88441, -77.35017, -77.35017,
  -77.88441, -77.88441, -77.35017, -77.35017,
  -77.35017, -77.35017, -76.81593, -76.81593,
  -77.35017, -77.35017, -76.81593, -76.81593,
  -77.35017, -77.35017, -76.81593, -76.81593,
  -77.35017, -77.35017, -76.81593, -76.81593,
  -77.35017, -77.35017, -76.81593, -76.81593,
  -77.35017, -77.35017, -76.81593, -76.81593,
  -77.35017, -77.35017, -76.81593, -76.81593,
  -77.35017, -77.35017, -76.81593, -76.81593,
  -77.35017, -77.35017, -76.81593, -76.81593,
  -77.35017, -77.35017, -76.81593, -76.81593,
  -77.35017, -77.35017, -76.81593, -76.81593,
  -77.35017, -77.35017, -76.81593, -76.81593,
  -77.35017, -77.35017, -76.81593, -76.81593,
  -77.35017, -77.35017, -76.81593, -76.81593,
  -77.35017, -77.35017, -76.81593, -76.81593,
  -77.35017, -77.35017, -76.81593, -76.81593,
  -77.35017, -77.35017, -76.81593, -76.81593,
  -77.35017, -77.35017, -76.81593, -76.81593,
  -77.35017, -77.35017, -76.81593, -76.81593,
  -77.35017, -77.35017, -76.81593, -76.81593,
  -76.81593, -76.81593, -76.28169, -76.28169,
  -76.81593, -76.81593, -76.28169, -76.28169,
  -76.81593, -76.81593, -76.28169, -76.28169,
  -76.81593, -76.81593, -76.28169, -76.28169,
  -76.81593, -76.81593, -76.28169, -76.28169,
  -76.81593, -76.81593, -76.28169, -76.28169,
  -76.81593, -76.81593, -76.28169, -76.28169,
  -76.81593, -76.81593, -76.28169, -76.28169,
  -76.81593, -76.81593, -76.28169, -76.28169,
  -76.81593, -76.81593, -76.28169, -76.28169,
  -76.81593, -76.81593, -76.28169, -76.28169,
  -76.81593, -76.81593, -76.28169, -76.28169,
  -76.81593, -76.81593, -76.28169, -76.28169,
  -76.81593, -76.81593, -76.28169, -76.28169,
  -76.81593, -76.81593, -76.28169, -76.28169,
  -76.81593, -76.81593, -76.28169, -76.28169,
  -76.81593, -76.81593, -76.28169, -76.28169,
  -76.81593, -76.81593, -76.28169, -76.28169,
  -76.81593, -76.81593, -76.28169, -76.28169,
  -76.81593, -76.81593, -76.28169, -76.28169,
  -76.28169, -76.28169, -75.74745, -75.74745,
  -76.28169, -76.28169, -75.74745, -75.74745,
  -76.28169, -76.28169, -75.74745, -75.74745,
  -76.28169, -76.28169, -75.74745, -75.74745,
  -76.28169, -76.28169, -75.74745, -75.74745,
  -76.28169, -76.28169, -75.74745, -75.74745,
  -76.28169, -76.28169, -75.74745, -75.74745,
  -76.28169, -76.28169, -75.74745, -75.74745,
  -76.28169, -76.28169, -75.74745, -75.74745,
  -76.28169, -76.28169, -75.74745, -75.74745,
  -76.28169, -76.28169, -75.74745, -75.74745,
  -76.28169, -76.28169, -75.74745, -75.74745,
  -76.28169, -76.28169, -75.74745, -75.74745,
  -76.28169, -76.28169, -75.74745, -75.74745,
  -76.28169, -76.28169, -75.74745, -75.74745,
  -76.28169, -76.28169, -75.74745, -75.74745,
  -76.28169, -76.28169, -75.74745, -75.74745,
  -76.28169, -76.28169, -75.74745, -75.74745,
  -76.28169, -76.28169, -75.74745, -75.74745,
  -76.28169, -76.28169, -75.74745, -75.74745,
  -75.74745, -75.74745, -75.21322, -75.21322,
  -75.74745, -75.74745, -75.21322, -75.21322,
  -75.74745, -75.74745, -75.21322, -75.21322,
  -75.74745, -75.74745, -75.21322, -75.21322,
  -75.74745, -75.74745, -75.21322, -75.21322,
  -75.74745, -75.74745, -75.21322, -75.21322,
  -75.74745, -75.74745, -75.21322, -75.21322,
  -75.74745, -75.74745, -75.21322, -75.21322,
  -75.74745, -75.74745, -75.21322, -75.21322,
  -75.74745, -75.74745, -75.21322, -75.21322,
  -75.74745, -75.74745, -75.21322, -75.21322,
  -75.74745, -75.74745, -75.21322, -75.21322,
  -75.74745, -75.74745, -75.21322, -75.21322,
  -75.74745, -75.74745, -75.21322, -75.21322,
  -75.74745, -75.74745, -75.21322, -75.21322,
  -75.74745, -75.74745, -75.21322, -75.21322,
  -75.74745, -75.74745, -75.21322, -75.21322,
  -75.74745, -75.74745, -75.21322, -75.21322,
  -75.74745, -75.74745, -75.21322, -75.21322,
  -75.74745, -75.74745, -75.21322, -75.21322,
  -75.21322, -75.21322, -74.67898, -74.67898,
  -75.21322, -75.21322, -74.67898, -74.67898,
  -75.21322, -75.21322, -74.67898, -74.67898,
  -75.21322, -75.21322, -74.67898, -74.67898,
  -75.21322, -75.21322, -74.67898, -74.67898,
  -75.21322, -75.21322, -74.67898, -74.67898,
  -75.21322, -75.21322, -74.67898, -74.67898,
  -75.21322, -75.21322, -74.67898, -74.67898,
  -75.21322, -75.21322, -74.67898, -74.67898,
  -75.21322, -75.21322, -74.67898, -74.67898,
  -75.21322, -75.21322, -74.67898, -74.67898,
  -75.21322, -75.21322, -74.67898, -74.67898,
  -75.21322, -75.21322, -74.67898, -74.67898,
  -75.21322, -75.21322, -74.67898, -74.67898,
  -75.21322, -75.21322, -74.67898, -74.67898,
  -75.21322, -75.21322, -74.67898, -74.67898,
  -75.21322, -75.21322, -74.67898, -74.67898,
  -75.21322, -75.21322, -74.67898, -74.67898,
  -75.21322, -75.21322, -74.67898, -74.67898,
  -75.21322, -75.21322, -74.67898, -74.67898,
  -74.67898, -74.67898, -74.14474, -74.14474,
  -74.67898, -74.67898, -74.14474, -74.14474,
  -74.67898, -74.67898, -74.14474, -74.14474,
  -74.67898, -74.67898, -74.14474, -74.14474,
  -74.67898, -74.67898, -74.14474, -74.14474,
  -74.67898, -74.67898, -74.14474, -74.14474,
  -74.67898, -74.67898, -74.14474, -74.14474,
  -74.67898, -74.67898, -74.14474, -74.14474,
  -74.67898, -74.67898, -74.14474, -74.14474,
  -74.67898, -74.67898, -74.14474, -74.14474,
  -74.67898, -74.67898, -74.14474, -74.14474,
  -74.67898, -74.67898, -74.14474, -74.14474,
  -74.67898, -74.67898, -74.14474, -74.14474,
  -74.67898, -74.67898, -74.14474, -74.14474,
  -74.67898, -74.67898, -74.14474, -74.14474,
  -74.67898, -74.67898, -74.14474, -74.14474,
  -74.67898, -74.67898, -74.14474, -74.14474,
  -74.67898, -74.67898, -74.14474, -74.14474,
  -74.67898, -74.67898, -74.14474, -74.14474,
  -74.67898, -74.67898, -74.14474, -74.14474,
  -74.14474, -74.14474, -73.6105, -73.6105,
  -74.14474, -74.14474, -73.6105, -73.6105,
  -74.14474, -74.14474, -73.6105, -73.6105,
  -74.14474, -74.14474, -73.6105, -73.6105,
  -74.14474, -74.14474, -73.6105, -73.6105,
  -74.14474, -74.14474, -73.6105, -73.6105,
  -74.14474, -74.14474, -73.6105, -73.6105,
  -74.14474, -74.14474, -73.6105, -73.6105,
  -74.14474, -74.14474, -73.6105, -73.6105,
  -74.14474, -74.14474, -73.6105, -73.6105,
  -74.14474, -74.14474, -73.6105, -73.6105,
  -74.14474, -74.14474, -73.6105, -73.6105,
  -74.14474, -74.14474, -73.6105, -73.6105,
  -74.14474, -74.14474, -73.6105, -73.6105,
  -74.14474, -74.14474, -73.6105, -73.6105,
  -74.14474, -74.14474, -73.6105, -73.6105,
  -74.14474, -74.14474, -73.6105, -73.6105,
  -74.14474, -74.14474, -73.6105, -73.6105,
  -74.14474, -74.14474, -73.6105, -73.6105,
  -74.14474, -74.14474, -73.6105, -73.6105,
  -73.6105, -73.6105, -73.07626, -73.07626,
  -73.6105, -73.6105, -73.07626, -73.07626,
  -73.6105, -73.6105, -73.07626, -73.07626,
  -73.6105, -73.6105, -73.07626, -73.07626,
  -73.6105, -73.6105, -73.07626, -73.07626,
  -73.6105, -73.6105, -73.07626, -73.07626,
  -73.6105, -73.6105, -73.07626, -73.07626,
  -73.6105, -73.6105, -73.07626, -73.07626,
  -73.6105, -73.6105, -73.07626, -73.07626,
  -73.6105, -73.6105, -73.07626, -73.07626,
  -73.6105, -73.6105, -73.07626, -73.07626,
  -73.6105, -73.6105, -73.07626, -73.07626,
  -73.6105, -73.6105, -73.07626, -73.07626,
  -73.6105, -73.6105, -73.07626, -73.07626,
  -73.6105, -73.6105, -73.07626, -73.07626,
  -73.6105, -73.6105, -73.07626, -73.07626,
  -73.6105, -73.6105, -73.07626, -73.07626,
  -73.6105, -73.6105, -73.07626, -73.07626,
  -73.6105, -73.6105, -73.07626, -73.07626,
  -73.6105, -73.6105, -73.07626, -73.07626,
  -73.07626, -73.07626, -72.54202, -72.54202,
  -73.07626, -73.07626, -72.54202, -72.54202,
  -73.07626, -73.07626, -72.54202, -72.54202,
  -73.07626, -73.07626, -72.54202, -72.54202,
  -73.07626, -73.07626, -72.54202, -72.54202,
  -73.07626, -73.07626, -72.54202, -72.54202,
  -73.07626, -73.07626, -72.54202, -72.54202,
  -73.07626, -73.07626, -72.54202, -72.54202,
  -73.07626, -73.07626, -72.54202, -72.54202,
  -73.07626, -73.07626, -72.54202, -72.54202,
  -73.07626, -73.07626, -72.54202, -72.54202,
  -73.07626, -73.07626, -72.54202, -72.54202,
  -73.07626, -73.07626, -72.54202, -72.54202,
  -73.07626, -73.07626, -72.54202, -72.54202,
  -73.07626, -73.07626, -72.54202, -72.54202,
  -73.07626, -73.07626, -72.54202, -72.54202,
  -73.07626, -73.07626, -72.54202, -72.54202,
  -73.07626, -73.07626, -72.54202, -72.54202,
  -73.07626, -73.07626, -72.54202, -72.54202,
  -73.07626, -73.07626, -72.54202, -72.54202,
  -72.54202, -72.54202, -72.00777, -72.00777,
  -72.54202, -72.54202, -72.00777, -72.00777,
  -72.54202, -72.54202, -72.00777, -72.00777,
  -72.54202, -72.54202, -72.00777, -72.00777,
  -72.54202, -72.54202, -72.00777, -72.00777,
  -72.54202, -72.54202, -72.00777, -72.00777,
  -72.54202, -72.54202, -72.00777, -72.00777,
  -72.54202, -72.54202, -72.00777, -72.00777,
  -72.54202, -72.54202, -72.00777, -72.00777,
  -72.54202, -72.54202, -72.00777, -72.00777,
  -72.54202, -72.54202, -72.00777, -72.00777,
  -72.54202, -72.54202, -72.00777, -72.00777,
  -72.54202, -72.54202, -72.00777, -72.00777,
  -72.54202, -72.54202, -72.00777, -72.00777,
  -72.54202, -72.54202, -72.00777, -72.00777,
  -72.54202, -72.54202, -72.00777, -72.00777,
  -72.54202, -72.54202, -72.00777, -72.00777,
  -72.54202, -72.54202, -72.00777, -72.00777,
  -72.54202, -72.54202, -72.00777, -72.00777,
  -72.54202, -72.54202, -72.00777, -72.00777,
  -72.00777, -72.00777, -71.47353, -71.47353,
  -72.00777, -72.00777, -71.47353, -71.47353,
  -72.00777, -72.00777, -71.47353, -71.47353,
  -72.00777, -72.00777, -71.47353, -71.47353,
  -72.00777, -72.00777, -71.47353, -71.47353,
  -72.00777, -72.00777, -71.47353, -71.47353,
  -72.00777, -72.00777, -71.47353, -71.47353,
  -72.00777, -72.00777, -71.47353, -71.47353,
  -72.00777, -72.00777, -71.47353, -71.47353,
  -72.00777, -72.00777, -71.47353, -71.47353,
  -72.00777, -72.00777, -71.47353, -71.47353,
  -72.00777, -72.00777, -71.47353, -71.47353,
  -72.00777, -72.00777, -71.47353, -71.47353,
  -72.00777, -72.00777, -71.47353, -71.47353,
  -72.00777, -72.00777, -71.47353, -71.47353,
  -72.00777, -72.00777, -71.47353, -71.47353,
  -72.00777, -72.00777, -71.47353, -71.47353,
  -72.00777, -72.00777, -71.47353, -71.47353,
  -72.00777, -72.00777, -71.47353, -71.47353,
  -72.00777, -72.00777, -71.47353, -71.47353,
  -71.47353, -71.47353, -70.93929, -70.93929,
  -71.47353, -71.47353, -70.93929, -70.93929,
  -71.47353, -71.47353, -70.93929, -70.93929,
  -71.47353, -71.47353, -70.93929, -70.93929,
  -71.47353, -71.47353, -70.93929, -70.93929,
  -71.47353, -71.47353, -70.93929, -70.93929,
  -71.47353, -71.47353, -70.93929, -70.93929,
  -71.47353, -71.47353, -70.93929, -70.93929,
  -71.47353, -71.47353, -70.93929, -70.93929,
  -71.47353, -71.47353, -70.93929, -70.93929,
  -71.47353, -71.47353, -70.93929, -70.93929,
  -71.47353, -71.47353, -70.93929, -70.93929,
  -71.47353, -71.47353, -70.93929, -70.93929,
  -71.47353, -71.47353, -70.93929, -70.93929,
  -71.47353, -71.47353, -70.93929, -70.93929,
  -71.47353, -71.47353, -70.93929, -70.93929,
  -71.47353, -71.47353, -70.93929, -70.93929,
  -71.47353, -71.47353, -70.93929, -70.93929,
  -71.47353, -71.47353, -70.93929, -70.93929,
  -71.47353, -71.47353, -70.93929, -70.93929,
  -70.93929, -70.93929, -70.40505, -70.40505,
  -70.93929, -70.93929, -70.40505, -70.40505,
  -70.93929, -70.93929, -70.40505, -70.40505,
  -70.93929, -70.93929, -70.40505, -70.40505,
  -70.93929, -70.93929, -70.40505, -70.40505,
  -70.93929, -70.93929, -70.40505, -70.40505,
  -70.93929, -70.93929, -70.40505, -70.40505,
  -70.93929, -70.93929, -70.40505, -70.40505,
  -70.93929, -70.93929, -70.40505, -70.40505,
  -70.93929, -70.93929, -70.40505, -70.40505,
  -70.93929, -70.93929, -70.40505, -70.40505,
  -70.93929, -70.93929, -70.40505, -70.40505,
  -70.93929, -70.93929, -70.40505, -70.40505,
  -70.93929, -70.93929, -70.40505, -70.40505,
  -70.93929, -70.93929, -70.40505, -70.40505,
  -70.93929, -70.93929, -70.40505, -70.40505,
  -70.93929, -70.93929, -70.40505, -70.40505,
  -70.93929, -70.93929, -70.40505, -70.40505,
  -70.93929, -70.93929, -70.40505, -70.40505,
  -70.93929, -70.93929, -70.40505, -70.40505,
  -70.40505, -70.40505, -69.87081, -69.87081,
  -70.40505, -70.40505, -69.87081, -69.87081,
  -70.40505, -70.40505, -69.87081, -69.87081,
  -70.40505, -70.40505, -69.87081, -69.87081,
  -70.40505, -70.40505, -69.87081, -69.87081,
  -70.40505, -70.40505, -69.87081, -69.87081,
  -70.40505, -70.40505, -69.87081, -69.87081,
  -70.40505, -70.40505, -69.87081, -69.87081,
  -70.40505, -70.40505, -69.87081, -69.87081,
  -70.40505, -70.40505, -69.87081, -69.87081,
  -70.40505, -70.40505, -69.87081, -69.87081,
  -70.40505, -70.40505, -69.87081, -69.87081,
  -70.40505, -70.40505, -69.87081, -69.87081,
  -70.40505, -70.40505, -69.87081, -69.87081,
  -70.40505, -70.40505, -69.87081, -69.87081,
  -70.40505, -70.40505, -69.87081, -69.87081,
  -70.40505, -70.40505, -69.87081, -69.87081,
  -70.40505, -70.40505, -69.87081, -69.87081,
  -70.40505, -70.40505, -69.87081, -69.87081,
  -70.40505, -70.40505, -69.87081, -69.87081,
  -69.87081, -69.87081, -69.33658, -69.33658,
  -69.87081, -69.87081, -69.33658, -69.33658,
  -69.87081, -69.87081, -69.33658, -69.33658,
  -69.87081, -69.87081, -69.33658, -69.33658,
  -69.87081, -69.87081, -69.33658, -69.33658,
  -69.87081, -69.87081, -69.33658, -69.33658,
  -69.87081, -69.87081, -69.33658, -69.33658,
  -69.87081, -69.87081, -69.33658, -69.33658,
  -69.87081, -69.87081, -69.33658, -69.33658,
  -69.87081, -69.87081, -69.33658, -69.33658,
  -69.87081, -69.87081, -69.33658, -69.33658,
  -69.87081, -69.87081, -69.33658, -69.33658,
  -69.87081, -69.87081, -69.33658, -69.33658,
  -69.87081, -69.87081, -69.33658, -69.33658,
  -69.87081, -69.87081, -69.33658, -69.33658,
  -69.87081, -69.87081, -69.33658, -69.33658,
  -69.87081, -69.87081, -69.33658, -69.33658,
  -69.87081, -69.87081, -69.33658, -69.33658,
  -69.87081, -69.87081, -69.33658, -69.33658,
  -69.87081, -69.87081, -69.33658, -69.33658,
  -69.33658, -69.33658, -68.80234, -68.80234,
  -69.33658, -69.33658, -68.80234, -68.80234,
  -69.33658, -69.33658, -68.80234, -68.80234,
  -69.33658, -69.33658, -68.80234, -68.80234,
  -69.33658, -69.33658, -68.80234, -68.80234,
  -69.33658, -69.33658, -68.80234, -68.80234,
  -69.33658, -69.33658, -68.80234, -68.80234,
  -69.33658, -69.33658, -68.80234, -68.80234,
  -69.33658, -69.33658, -68.80234, -68.80234,
  -69.33658, -69.33658, -68.80234, -68.80234,
  -69.33658, -69.33658, -68.80234, -68.80234,
  -69.33658, -69.33658, -68.80234, -68.80234,
  -69.33658, -69.33658, -68.80234, -68.80234,
  -69.33658, -69.33658, -68.80234, -68.80234,
  -69.33658, -69.33658, -68.80234, -68.80234,
  -69.33658, -69.33658, -68.80234, -68.80234,
  -69.33658, -69.33658, -68.80234, -68.80234,
  -69.33658, -69.33658, -68.80234, -68.80234,
  -69.33658, -69.33658, -68.80234, -68.80234,
  -69.33658, -69.33658, -68.80234, -68.80234 ;

 time = 18265.5, 18295, 18324.5, 18355 ;

 time_bnds =
  18250, 18281,
  18281, 18309,
  18309, 18340,
  18340, 18370 ;

 sos =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  33.82447, 33.82838, 33.84248, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  33.78296, 33.81977, 33.83622, 33.82368, 33.8135, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  33.84562, 33.89261, 33.90436, 33.88008, 33.83152, 33.77747, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  33.97015, 33.99678, 34.00305, 33.96232, 33.90749, 33.85423, 33.79705, 
    33.79784, 33.82133, _, _, _, _, _, _, _, _, _, _, _,
  34.08921, 34.07589, 34.04143, 34.02342, 34.00305, 33.97094, 33.94039, 
    33.91298, 33.87773, 33.83543, 33.83935, _, _, _, _, _, _, _, _, _,
  34.13307, 34.09313, 34.05318, 34.03673, 34.0195, 34.00227, 33.97485, 
    33.95449, 33.91768, 33.87146, 33.84718, 33.79314, _, _, _, _, _, _, _, _,
  34.11662, 34.09156, 34.06415, 34.0383, 34.0195, 33.99287, 33.96624, 
    33.92629, 33.88869, 33.87146, 33.83935, 33.77434, 33.70855, _, _, _, _, 
    _, _, _,
  34.05553, 34.03673, 34.02811, 34.01558, 34.00227, 33.98347, 33.94744, 
    33.89261, 33.85501, 33.83543, 33.81977, 33.76886, 33.66703, _, _, _, _, 
    _, _, _,
  33.98738, 33.98269, 33.97799, 33.97015, 33.94822, 33.92551, 33.88321, 
    33.84483, 33.81037, 33.78531, 33.75163, 33.70228, 33.66233, 33.64354, _, 
    _, _, _, _, _,
  33.94666, 33.95527, 33.9584, 33.94587, 33.92081, 33.88791, 33.8558, 
    33.82212, 33.79157, 33.76886, 33.74536, 33.70776, 33.67408, 33.64119, 
    33.61847, 33.60751, 33.58322, _, _, _,
  33.92707, 33.94117, 33.94744, 33.94431, 33.92629, 33.89966, 33.86363, 
    33.83073, 33.79705, 33.77356, 33.75084, 33.72813, 33.70228, 33.66312, 
    33.62082, 33.59262, 33.56756, 33.53936, _, _,
  33.90123, 33.92159, 33.93491, 33.93099, 33.91298, 33.89418, 33.86676, 
    33.84483, 33.81977, 33.7994, 33.78609, 33.76807, 33.74771, 33.72108, 
    33.69836, 33.67095, 33.63022, 33.59889, 33.59262, 33.58479,
  33.86285, 33.8793, 33.89104, 33.89574, 33.88869, 33.8793, 33.86128, 
    33.84875, 33.837, 33.82682, 33.81507, 33.81115, 33.81742, 33.81585, 
    33.80254, 33.77434, 33.74066, 33.71325, 33.70855, 33.69993,
  33.81429, 33.83857, 33.85736, 33.86598, 33.86441, 33.86206, 33.85815, 
    33.85893, 33.85658, 33.85423, 33.85032, 33.85188, 33.85501, 33.85893, 
    33.85658, 33.84797, 33.83935, 33.84013, 33.84797, 33.84327,
  33.75163, 33.77512, 33.80097, 33.82682, 33.84562, 33.85345, 33.85658, 
    33.86128, 33.86598, 33.8699, 33.86755, 33.8652, 33.86911, 33.88008, 
    33.88869, 33.89418, 33.89653, 33.90123, 33.90906, 33.91376,
  33.69915, 33.72578, 33.75476, 33.77747, 33.79784, 33.8135, 33.82525, 
    33.83857, 33.84875, 33.85423, 33.85423, 33.85345, 33.85423, 33.86911, 
    33.88791, 33.90279, 33.91611, 33.93099, 33.94196, 33.94744,
  33.68818, 33.68505, 33.69053, 33.71638, 33.74536, 33.76181, 33.76886, 
    33.77356, 33.77591, 33.77669, 33.77982, 33.78531, 33.7947, 33.81272, 
    33.83465, 33.85501, 33.87616, 33.90123, 33.92707, 33.94822,
  33.72343, 33.70463, 33.68427, 33.67487, 33.67957, 33.68975, 33.69601, 
    33.69836, 33.69131, 33.68113, 33.67252, 33.67095, 33.6733, 33.68975, 
    33.71168, 33.73518, 33.75867, 33.78844, 33.82525, 33.86363,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  33.87363, 33.87912, 33.88225, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  33.86031, 33.88382, 33.88695, 33.87285, 33.86266, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  33.96216, 33.97626, 33.97548, 33.94571, 33.89557, 33.83211, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  33.99506, 34.01073, 34.01308, 33.98723, 33.95041, 33.90654, 33.85483, 
    33.85483, 33.85796, _, _, _, _, _, _, _, _, _, _, _,
  34.0452, 34.0452, 34.02326, 34.01308, 34.0029, 33.98566, 33.96216, 
    33.94414, 33.90575, 33.85405, 33.83446, _, _, _, _, _, _, _, _, _,
  34.1016, 34.06244, 34.02718, 34.01308, 34.00211, 33.99506, 33.98018, 
    33.96373, 33.93004, 33.88773, 33.84386, 33.79294, _, _, _, _, _, _, _, _,
  34.10395, 34.08358, 34.04755, 34.01464, 33.98958, 33.96999, 33.95275, 
    33.93317, 33.92455, 33.89557, 33.84465, 33.77649, 33.71852, _, _, _, _, 
    _, _, _,
  34.05303, 34.02561, 34.0029, 33.98331, 33.96686, 33.95275, 33.91907, 
    33.87833, 33.85561, 33.83211, 33.80626, 33.78041, 33.72557, _, _, _, _, 
    _, _, _,
  33.96999, 33.96294, 33.95197, 33.93317, 33.90967, 33.88773, 33.85405, 
    33.82193, 33.79843, 33.77884, 33.74124, 33.70834, 33.68718, 33.64175, _, 
    _, _, _, _, _,
  33.93082, 33.93866, 33.93317, 33.90967, 33.87912, 33.84621, 33.82036, 
    33.79137, 33.76631, 33.74751, 33.72322, 33.69423, 33.67073, 33.64331, 
    33.61589, 33.59709, 33.57751, _, _, _,
  33.91202, 33.92455, 33.92455, 33.90497, 33.87598, 33.84386, 33.81644, 
    33.78981, 33.76631, 33.74672, 33.72087, 33.6958, 33.66838, 33.64018, 
    33.60728, 33.57829, 33.55714, 33.52815, _, _,
  33.89322, 33.90732, 33.9081, 33.89322, 33.87207, 33.84465, 33.82114, 
    33.80234, 33.78746, 33.77649, 33.76082, 33.73732, 33.71304, 33.68562, 
    33.65115, 33.61354, 33.57751, 33.55635, 33.55009, 33.5493,
  33.86266, 33.87442, 33.87755, 33.86893, 33.85483, 33.83916, 33.82584, 
    33.81801, 33.81096, 33.80626, 33.80313, 33.79921, 33.78981, 33.77101, 
    33.7381, 33.70128, 33.66838, 33.65036, 33.65193, 33.64331,
  33.82349, 33.83916, 33.84621, 33.84465, 33.83995, 33.83525, 33.83368, 
    33.8329, 33.83133, 33.83055, 33.8329, 33.8376, 33.84073, 33.83446, 
    33.81958, 33.80156, 33.78667, 33.77962, 33.78041, 33.77414,
  33.76866, 33.78589, 33.80234, 33.81331, 33.81958, 33.82428, 33.82898, 
    33.83211, 33.8329, 33.83211, 33.83133, 33.83446, 33.84386, 33.85405, 
    33.8611, 33.86345, 33.86345, 33.86345, 33.86502, 33.86188,
  33.71069, 33.73027, 33.75299, 33.77022, 33.78511, 33.79686, 33.80548, 
    33.80704, 33.80548, 33.79843, 33.79216, 33.79216, 33.80313, 33.82428, 
    33.84778, 33.86658, 33.87912, 33.89008, 33.89714, 33.89949,
  33.66211, 33.67387, 33.69423, 33.71695, 33.73654, 33.74751, 33.74986, 
    33.74359, 33.73262, 33.71225, 33.69658, 33.69267, 33.70363, 33.72713, 
    33.75455, 33.78119, 33.80469, 33.83133, 33.8564, 33.8752,
  33.6535, 33.64331, 33.65115, 33.67073, 33.69188, 33.69972, 33.69345, 
    33.67387, 33.64331, 33.61041, 33.57907, 33.5634, 33.56419, 33.57594, 
    33.59474, 33.61903, 33.65193, 33.69501, 33.74359, 33.77806,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  33.88458, 33.8838, 33.8838, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  33.87753, 33.89241, 33.89241, 33.87283, 33.86265, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  33.99188, 33.99345, 33.97935, 33.94489, 33.89633, 33.84151, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  34.06707, 34.05062, 34.02791, 33.99345, 33.94724, 33.9026, 33.85091, 
    33.84621, 33.84229, _, _, _, _, _, _, _, _, _, _, _,
  34.12816, 34.10937, 34.06316, 34.03339, 34.01068, 33.9864, 33.96291, 
    33.94411, 33.8979, 33.83524, 33.81253, _, _, _, _, _, _, _, _, _,
  34.18534, 34.13599, 34.08822, 34.05376, 34.02791, 34.01146, 33.99502, 
    33.97309, 33.93941, 33.90181, 33.85482, 33.8, _, _, _, _, _, _, _, _,
  34.1916, 34.16576, 34.11485, 34.06864, 34.02791, 33.99815, 33.97465, 
    33.95977, 33.95351, 33.93079, 33.87127, 33.80078, 33.73342, _, _, _, _, 
    _, _, _,
  34.15636, 34.12738, 34.08665, 34.05689, 34.02399, 33.9864, 33.93941, 
    33.89633, 33.87362, 33.85874, 33.82898, 33.81253, 33.7718, _, _, _, _, _, 
    _, _,
  34.07099, 34.05532, 34.02869, 34.00128, 33.97622, 33.94254, 33.89241, 
    33.85169, 33.81801, 33.80156, 33.78355, 33.77102, 33.74439, 33.69975, _, 
    _, _, _, _, _,
  34.02634, 34.01773, 33.99815, 33.96604, 33.93393, 33.90103, 33.87048, 
    33.83759, 33.8047, 33.78355, 33.76788, 33.75613, 33.74125, 33.71463, 
    33.67703, 33.6504, 33.62769, _, _, _,
  34.01303, 34.00285, 33.98249, 33.95272, 33.92296, 33.89555, 33.87127, 
    33.84542, 33.81723, 33.79216, 33.76945, 33.75457, 33.74125, 33.72481, 
    33.70366, 33.68095, 33.6551, 33.62534, _, _,
  33.99345, 33.9864, 33.96917, 33.94567, 33.92296, 33.90025, 33.88067, 
    33.86344, 33.84699, 33.82976, 33.80939, 33.78668, 33.76867, 33.74909, 
    33.73107, 33.70993, 33.69191, 33.67311, 33.66058, 33.66842,
  33.96682, 33.96212, 33.94881, 33.93314, 33.91748, 33.90338, 33.89241, 
    33.8838, 33.87597, 33.86735, 33.85795, 33.84542, 33.82898, 33.80704, 
    33.78511, 33.76318, 33.75144, 33.74439, 33.74752, 33.76005,
  33.93393, 33.93158, 33.92688, 33.91748, 33.91043, 33.90651, 33.90338, 
    33.89946, 33.89398, 33.89006, 33.88771, 33.88693, 33.88223, 33.87127, 
    33.8556, 33.84072, 33.83289, 33.83289, 33.84307, 33.85169,
  33.8885, 33.89241, 33.89711, 33.89476, 33.89398, 33.8932, 33.89633, 
    33.89476, 33.89241, 33.88928, 33.88693, 33.8885, 33.89241, 33.89633, 
    33.89711, 33.89476, 33.8932, 33.8932, 33.8979, 33.90025,
  33.83916, 33.84621, 33.85795, 33.86265, 33.86735, 33.87048, 33.87127, 
    33.86813, 33.86265, 33.85482, 33.84856, 33.84934, 33.8603, 33.87675, 
    33.89006, 33.90103, 33.9073, 33.91278, 33.91669, 33.91904,
  33.79921, 33.80626, 33.81879, 33.82976, 33.83759, 33.83916, 33.83211, 
    33.82114, 33.80704, 33.79373, 33.78355, 33.78198, 33.79373, 33.81253, 
    33.83211, 33.85091, 33.86735, 33.87988, 33.89241, 33.90103,
  33.7859, 33.78746, 33.80078, 33.81879, 33.82819, 33.82506, 33.81174, 
    33.7906, 33.76632, 33.74595, 33.73421, 33.73029, 33.73734, 33.75144, 
    33.76867, 33.78746, 33.81174, 33.83446, 33.85325, 33.86422,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  33.83966, 33.8154, 33.81853, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  33.79349, 33.82792, 33.84357, 33.82166, 33.81931, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  33.93357, 33.93357, 33.94765, 33.91244, 33.86861, 33.80523, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  34.09321, 34.10651, 34.07834, 34.04, 33.98209, 33.91792, 33.87409, 
    33.85609, 33.84748, _, _, _, _, _, _, _, _, _, _, _,
  34.2286, 34.19886, 34.14721, 34.10495, 34.07521, 34.0533, 34.02513, 
    34.00087, 33.94609, 33.88427, 33.84357, _, _, _, _, _, _, _, _, _,
  34.2646, 34.22546, 34.18164, 34.14643, 34.11434, 34.09321, 34.07443, 
    34.0533, 34.02435, 33.98913, 33.93904, 33.87879, _, _, _, _, _, _, _, _,
  34.24347, 34.23642, 34.20042, 34.15425, 34.10886, 34.07756, 34.05487, 
    34.04156, 34.03608, 34.02356, 33.98365, 33.90931, 33.82401, _, _, _, _, 
    _, _, _,
  34.22781, 34.2059, 34.16677, 34.13547, 34.09947, 34.05643, 34.01261, 
    33.97504, 33.95391, 33.94218, 33.92809, 33.91557, 33.86314, _, _, _, _, 
    _, _, _,
  34.16051, 34.13704, 34.10808, 34.076, 34.04704, 34.00478, 33.95705, 
    33.9187, 33.88896, 33.87487, 33.87018, 33.86157, 33.82479, 33.76923, _, 
    _, _, _, _, _,
  34.11043, 34.0893, 34.06269, 34.02904, 33.99617, 33.96174, 33.93044, 
    33.89835, 33.86783, 33.85218, 33.84357, 33.83653, 33.82088, 33.78175, 
    33.72775, 33.68784, 33.66906, _, _, _,
  34.09321, 34.0666, 34.03765, 34.00713, 33.97818, 33.95078, 33.92731, 
    33.90226, 33.87644, 33.85688, 33.84044, 33.83262, 33.82088, 33.79975, 
    33.77079, 33.74497, 33.72149, 33.68393, _, _,
  34.07912, 34.05408, 34.02748, 34.00165, 33.97896, 33.95705, 33.93826, 
    33.92183, 33.90383, 33.88818, 33.87096, 33.85296, 33.8381, 33.82479, 
    33.81384, 33.79897, 33.77549, 33.74419, 33.72149, 33.73401,
  34.06034, 34.04, 34.01887, 34.00009, 33.98365, 33.96957, 33.95626, 33.9453, 
    33.93357, 33.92418, 33.91401, 33.89992, 33.88427, 33.86783, 33.85374, 
    33.84044, 33.83105, 33.81931, 33.8107, 33.8334,
  34.04078, 34.02591, 34.01417, 34.00009, 33.9907, 33.98365, 33.97583, 
    33.96487, 33.95548, 33.95, 33.94609, 33.94139, 33.93279, 33.9187, 
    33.9054, 33.89679, 33.88974, 33.89366, 33.90305, 33.91635,
  34.01495, 34.00791, 34.00322, 33.99617, 33.98913, 33.98365, 33.97896, 
    33.97113, 33.96487, 33.95783, 33.9547, 33.95313, 33.95235, 33.94844, 
    33.94452, 33.93826, 33.93435, 33.93435, 33.93904, 33.9453,
  33.98756, 33.986, 33.98522, 33.98522, 33.98287, 33.97896, 33.97191, 
    33.96409, 33.95783, 33.94922, 33.94374, 33.94374, 33.94922, 33.95391, 
    33.95705, 33.95626, 33.9547, 33.95548, 33.95626, 33.95626,
  33.96878, 33.97035, 33.97426, 33.97661, 33.97818, 33.97426, 33.96409, 
    33.95313, 33.94374, 33.93435, 33.92809, 33.92809, 33.93513, 33.94452, 
    33.95235, 33.95705, 33.96017, 33.96174, 33.96096, 33.95783,
  33.97426, 33.97818, 33.98522, 33.9907, 33.99226, 33.98678, 33.97583, 
    33.95861, 33.94139, 33.93044, 33.92731, 33.92887, 33.93513, 33.94452, 
    33.95391, 33.96409, 33.97035, 33.97191, 33.96957, 33.96565 ;
}
